magic
tech sky130B
magscale 1 2
timestamp 1662906990
<< obsli1 >>
rect 1104 2159 558808 497777
<< obsm1 >>
rect 1104 144 558808 499588
<< metal2 >>
rect 4894 499200 4950 500000
rect 9678 499200 9734 500000
rect 14462 499200 14518 500000
rect 19246 499200 19302 500000
rect 24030 499200 24086 500000
rect 28814 499200 28870 500000
rect 33598 499200 33654 500000
rect 38382 499200 38438 500000
rect 43166 499200 43222 500000
rect 47950 499200 48006 500000
rect 52734 499200 52790 500000
rect 57518 499200 57574 500000
rect 62302 499200 62358 500000
rect 67086 499200 67142 500000
rect 71870 499200 71926 500000
rect 76654 499200 76710 500000
rect 81438 499200 81494 500000
rect 86222 499200 86278 500000
rect 91006 499200 91062 500000
rect 95790 499200 95846 500000
rect 100574 499200 100630 500000
rect 105358 499200 105414 500000
rect 110142 499200 110198 500000
rect 114926 499200 114982 500000
rect 119710 499200 119766 500000
rect 124494 499200 124550 500000
rect 129278 499200 129334 500000
rect 134062 499200 134118 500000
rect 138846 499200 138902 500000
rect 143630 499200 143686 500000
rect 148414 499200 148470 500000
rect 153198 499200 153254 500000
rect 157982 499200 158038 500000
rect 162766 499200 162822 500000
rect 167550 499200 167606 500000
rect 172334 499200 172390 500000
rect 177118 499200 177174 500000
rect 181902 499200 181958 500000
rect 186686 499200 186742 500000
rect 191470 499200 191526 500000
rect 196254 499200 196310 500000
rect 201038 499200 201094 500000
rect 205822 499200 205878 500000
rect 210606 499200 210662 500000
rect 215390 499200 215446 500000
rect 220174 499200 220230 500000
rect 224958 499200 225014 500000
rect 229742 499200 229798 500000
rect 234526 499200 234582 500000
rect 239310 499200 239366 500000
rect 244094 499200 244150 500000
rect 248878 499200 248934 500000
rect 253662 499200 253718 500000
rect 258446 499200 258502 500000
rect 263230 499200 263286 500000
rect 268014 499200 268070 500000
rect 272798 499200 272854 500000
rect 277582 499200 277638 500000
rect 282366 499200 282422 500000
rect 287150 499200 287206 500000
rect 291934 499200 291990 500000
rect 296718 499200 296774 500000
rect 301502 499200 301558 500000
rect 306286 499200 306342 500000
rect 311070 499200 311126 500000
rect 315854 499200 315910 500000
rect 320638 499200 320694 500000
rect 325422 499200 325478 500000
rect 330206 499200 330262 500000
rect 334990 499200 335046 500000
rect 339774 499200 339830 500000
rect 344558 499200 344614 500000
rect 349342 499200 349398 500000
rect 354126 499200 354182 500000
rect 358910 499200 358966 500000
rect 363694 499200 363750 500000
rect 368478 499200 368534 500000
rect 373262 499200 373318 500000
rect 378046 499200 378102 500000
rect 382830 499200 382886 500000
rect 387614 499200 387670 500000
rect 392398 499200 392454 500000
rect 397182 499200 397238 500000
rect 401966 499200 402022 500000
rect 406750 499200 406806 500000
rect 411534 499200 411590 500000
rect 416318 499200 416374 500000
rect 421102 499200 421158 500000
rect 425886 499200 425942 500000
rect 430670 499200 430726 500000
rect 435454 499200 435510 500000
rect 440238 499200 440294 500000
rect 445022 499200 445078 500000
rect 449806 499200 449862 500000
rect 454590 499200 454646 500000
rect 459374 499200 459430 500000
rect 464158 499200 464214 500000
rect 468942 499200 468998 500000
rect 473726 499200 473782 500000
rect 478510 499200 478566 500000
rect 483294 499200 483350 500000
rect 488078 499200 488134 500000
rect 492862 499200 492918 500000
rect 497646 499200 497702 500000
rect 502430 499200 502486 500000
rect 507214 499200 507270 500000
rect 511998 499200 512054 500000
rect 516782 499200 516838 500000
rect 521566 499200 521622 500000
rect 526350 499200 526406 500000
rect 531134 499200 531190 500000
rect 535918 499200 535974 500000
rect 540702 499200 540758 500000
rect 545486 499200 545542 500000
rect 550270 499200 550326 500000
rect 555054 499200 555110 500000
rect 6090 0 6146 800
rect 7286 0 7342 800
rect 8482 0 8538 800
rect 9678 0 9734 800
rect 10874 0 10930 800
rect 12070 0 12126 800
rect 13266 0 13322 800
rect 14462 0 14518 800
rect 15658 0 15714 800
rect 16854 0 16910 800
rect 18050 0 18106 800
rect 19246 0 19302 800
rect 20442 0 20498 800
rect 21638 0 21694 800
rect 22834 0 22890 800
rect 24030 0 24086 800
rect 25226 0 25282 800
rect 26422 0 26478 800
rect 27618 0 27674 800
rect 28814 0 28870 800
rect 30010 0 30066 800
rect 31206 0 31262 800
rect 32402 0 32458 800
rect 33598 0 33654 800
rect 34794 0 34850 800
rect 35990 0 36046 800
rect 37186 0 37242 800
rect 38382 0 38438 800
rect 39578 0 39634 800
rect 40774 0 40830 800
rect 41970 0 42026 800
rect 43166 0 43222 800
rect 44362 0 44418 800
rect 45558 0 45614 800
rect 46754 0 46810 800
rect 47950 0 48006 800
rect 49146 0 49202 800
rect 50342 0 50398 800
rect 51538 0 51594 800
rect 52734 0 52790 800
rect 53930 0 53986 800
rect 55126 0 55182 800
rect 56322 0 56378 800
rect 57518 0 57574 800
rect 58714 0 58770 800
rect 59910 0 59966 800
rect 61106 0 61162 800
rect 62302 0 62358 800
rect 63498 0 63554 800
rect 64694 0 64750 800
rect 65890 0 65946 800
rect 67086 0 67142 800
rect 68282 0 68338 800
rect 69478 0 69534 800
rect 70674 0 70730 800
rect 71870 0 71926 800
rect 73066 0 73122 800
rect 74262 0 74318 800
rect 75458 0 75514 800
rect 76654 0 76710 800
rect 77850 0 77906 800
rect 79046 0 79102 800
rect 80242 0 80298 800
rect 81438 0 81494 800
rect 82634 0 82690 800
rect 83830 0 83886 800
rect 85026 0 85082 800
rect 86222 0 86278 800
rect 87418 0 87474 800
rect 88614 0 88670 800
rect 89810 0 89866 800
rect 91006 0 91062 800
rect 92202 0 92258 800
rect 93398 0 93454 800
rect 94594 0 94650 800
rect 95790 0 95846 800
rect 96986 0 97042 800
rect 98182 0 98238 800
rect 99378 0 99434 800
rect 100574 0 100630 800
rect 101770 0 101826 800
rect 102966 0 103022 800
rect 104162 0 104218 800
rect 105358 0 105414 800
rect 106554 0 106610 800
rect 107750 0 107806 800
rect 108946 0 109002 800
rect 110142 0 110198 800
rect 111338 0 111394 800
rect 112534 0 112590 800
rect 113730 0 113786 800
rect 114926 0 114982 800
rect 116122 0 116178 800
rect 117318 0 117374 800
rect 118514 0 118570 800
rect 119710 0 119766 800
rect 120906 0 120962 800
rect 122102 0 122158 800
rect 123298 0 123354 800
rect 124494 0 124550 800
rect 125690 0 125746 800
rect 126886 0 126942 800
rect 128082 0 128138 800
rect 129278 0 129334 800
rect 130474 0 130530 800
rect 131670 0 131726 800
rect 132866 0 132922 800
rect 134062 0 134118 800
rect 135258 0 135314 800
rect 136454 0 136510 800
rect 137650 0 137706 800
rect 138846 0 138902 800
rect 140042 0 140098 800
rect 141238 0 141294 800
rect 142434 0 142490 800
rect 143630 0 143686 800
rect 144826 0 144882 800
rect 146022 0 146078 800
rect 147218 0 147274 800
rect 148414 0 148470 800
rect 149610 0 149666 800
rect 150806 0 150862 800
rect 152002 0 152058 800
rect 153198 0 153254 800
rect 154394 0 154450 800
rect 155590 0 155646 800
rect 156786 0 156842 800
rect 157982 0 158038 800
rect 159178 0 159234 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162766 0 162822 800
rect 163962 0 164018 800
rect 165158 0 165214 800
rect 166354 0 166410 800
rect 167550 0 167606 800
rect 168746 0 168802 800
rect 169942 0 169998 800
rect 171138 0 171194 800
rect 172334 0 172390 800
rect 173530 0 173586 800
rect 174726 0 174782 800
rect 175922 0 175978 800
rect 177118 0 177174 800
rect 178314 0 178370 800
rect 179510 0 179566 800
rect 180706 0 180762 800
rect 181902 0 181958 800
rect 183098 0 183154 800
rect 184294 0 184350 800
rect 185490 0 185546 800
rect 186686 0 186742 800
rect 187882 0 187938 800
rect 189078 0 189134 800
rect 190274 0 190330 800
rect 191470 0 191526 800
rect 192666 0 192722 800
rect 193862 0 193918 800
rect 195058 0 195114 800
rect 196254 0 196310 800
rect 197450 0 197506 800
rect 198646 0 198702 800
rect 199842 0 199898 800
rect 201038 0 201094 800
rect 202234 0 202290 800
rect 203430 0 203486 800
rect 204626 0 204682 800
rect 205822 0 205878 800
rect 207018 0 207074 800
rect 208214 0 208270 800
rect 209410 0 209466 800
rect 210606 0 210662 800
rect 211802 0 211858 800
rect 212998 0 213054 800
rect 214194 0 214250 800
rect 215390 0 215446 800
rect 216586 0 216642 800
rect 217782 0 217838 800
rect 218978 0 219034 800
rect 220174 0 220230 800
rect 221370 0 221426 800
rect 222566 0 222622 800
rect 223762 0 223818 800
rect 224958 0 225014 800
rect 226154 0 226210 800
rect 227350 0 227406 800
rect 228546 0 228602 800
rect 229742 0 229798 800
rect 230938 0 230994 800
rect 232134 0 232190 800
rect 233330 0 233386 800
rect 234526 0 234582 800
rect 235722 0 235778 800
rect 236918 0 236974 800
rect 238114 0 238170 800
rect 239310 0 239366 800
rect 240506 0 240562 800
rect 241702 0 241758 800
rect 242898 0 242954 800
rect 244094 0 244150 800
rect 245290 0 245346 800
rect 246486 0 246542 800
rect 247682 0 247738 800
rect 248878 0 248934 800
rect 250074 0 250130 800
rect 251270 0 251326 800
rect 252466 0 252522 800
rect 253662 0 253718 800
rect 254858 0 254914 800
rect 256054 0 256110 800
rect 257250 0 257306 800
rect 258446 0 258502 800
rect 259642 0 259698 800
rect 260838 0 260894 800
rect 262034 0 262090 800
rect 263230 0 263286 800
rect 264426 0 264482 800
rect 265622 0 265678 800
rect 266818 0 266874 800
rect 268014 0 268070 800
rect 269210 0 269266 800
rect 270406 0 270462 800
rect 271602 0 271658 800
rect 272798 0 272854 800
rect 273994 0 274050 800
rect 275190 0 275246 800
rect 276386 0 276442 800
rect 277582 0 277638 800
rect 278778 0 278834 800
rect 279974 0 280030 800
rect 281170 0 281226 800
rect 282366 0 282422 800
rect 283562 0 283618 800
rect 284758 0 284814 800
rect 285954 0 286010 800
rect 287150 0 287206 800
rect 288346 0 288402 800
rect 289542 0 289598 800
rect 290738 0 290794 800
rect 291934 0 291990 800
rect 293130 0 293186 800
rect 294326 0 294382 800
rect 295522 0 295578 800
rect 296718 0 296774 800
rect 297914 0 297970 800
rect 299110 0 299166 800
rect 300306 0 300362 800
rect 301502 0 301558 800
rect 302698 0 302754 800
rect 303894 0 303950 800
rect 305090 0 305146 800
rect 306286 0 306342 800
rect 307482 0 307538 800
rect 308678 0 308734 800
rect 309874 0 309930 800
rect 311070 0 311126 800
rect 312266 0 312322 800
rect 313462 0 313518 800
rect 314658 0 314714 800
rect 315854 0 315910 800
rect 317050 0 317106 800
rect 318246 0 318302 800
rect 319442 0 319498 800
rect 320638 0 320694 800
rect 321834 0 321890 800
rect 323030 0 323086 800
rect 324226 0 324282 800
rect 325422 0 325478 800
rect 326618 0 326674 800
rect 327814 0 327870 800
rect 329010 0 329066 800
rect 330206 0 330262 800
rect 331402 0 331458 800
rect 332598 0 332654 800
rect 333794 0 333850 800
rect 334990 0 335046 800
rect 336186 0 336242 800
rect 337382 0 337438 800
rect 338578 0 338634 800
rect 339774 0 339830 800
rect 340970 0 341026 800
rect 342166 0 342222 800
rect 343362 0 343418 800
rect 344558 0 344614 800
rect 345754 0 345810 800
rect 346950 0 347006 800
rect 348146 0 348202 800
rect 349342 0 349398 800
rect 350538 0 350594 800
rect 351734 0 351790 800
rect 352930 0 352986 800
rect 354126 0 354182 800
rect 355322 0 355378 800
rect 356518 0 356574 800
rect 357714 0 357770 800
rect 358910 0 358966 800
rect 360106 0 360162 800
rect 361302 0 361358 800
rect 362498 0 362554 800
rect 363694 0 363750 800
rect 364890 0 364946 800
rect 366086 0 366142 800
rect 367282 0 367338 800
rect 368478 0 368534 800
rect 369674 0 369730 800
rect 370870 0 370926 800
rect 372066 0 372122 800
rect 373262 0 373318 800
rect 374458 0 374514 800
rect 375654 0 375710 800
rect 376850 0 376906 800
rect 378046 0 378102 800
rect 379242 0 379298 800
rect 380438 0 380494 800
rect 381634 0 381690 800
rect 382830 0 382886 800
rect 384026 0 384082 800
rect 385222 0 385278 800
rect 386418 0 386474 800
rect 387614 0 387670 800
rect 388810 0 388866 800
rect 390006 0 390062 800
rect 391202 0 391258 800
rect 392398 0 392454 800
rect 393594 0 393650 800
rect 394790 0 394846 800
rect 395986 0 396042 800
rect 397182 0 397238 800
rect 398378 0 398434 800
rect 399574 0 399630 800
rect 400770 0 400826 800
rect 401966 0 402022 800
rect 403162 0 403218 800
rect 404358 0 404414 800
rect 405554 0 405610 800
rect 406750 0 406806 800
rect 407946 0 408002 800
rect 409142 0 409198 800
rect 410338 0 410394 800
rect 411534 0 411590 800
rect 412730 0 412786 800
rect 413926 0 413982 800
rect 415122 0 415178 800
rect 416318 0 416374 800
rect 417514 0 417570 800
rect 418710 0 418766 800
rect 419906 0 419962 800
rect 421102 0 421158 800
rect 422298 0 422354 800
rect 423494 0 423550 800
rect 424690 0 424746 800
rect 425886 0 425942 800
rect 427082 0 427138 800
rect 428278 0 428334 800
rect 429474 0 429530 800
rect 430670 0 430726 800
rect 431866 0 431922 800
rect 433062 0 433118 800
rect 434258 0 434314 800
rect 435454 0 435510 800
rect 436650 0 436706 800
rect 437846 0 437902 800
rect 439042 0 439098 800
rect 440238 0 440294 800
rect 441434 0 441490 800
rect 442630 0 442686 800
rect 443826 0 443882 800
rect 445022 0 445078 800
rect 446218 0 446274 800
rect 447414 0 447470 800
rect 448610 0 448666 800
rect 449806 0 449862 800
rect 451002 0 451058 800
rect 452198 0 452254 800
rect 453394 0 453450 800
rect 454590 0 454646 800
rect 455786 0 455842 800
rect 456982 0 457038 800
rect 458178 0 458234 800
rect 459374 0 459430 800
rect 460570 0 460626 800
rect 461766 0 461822 800
rect 462962 0 463018 800
rect 464158 0 464214 800
rect 465354 0 465410 800
rect 466550 0 466606 800
rect 467746 0 467802 800
rect 468942 0 468998 800
rect 470138 0 470194 800
rect 471334 0 471390 800
rect 472530 0 472586 800
rect 473726 0 473782 800
rect 474922 0 474978 800
rect 476118 0 476174 800
rect 477314 0 477370 800
rect 478510 0 478566 800
rect 479706 0 479762 800
rect 480902 0 480958 800
rect 482098 0 482154 800
rect 483294 0 483350 800
rect 484490 0 484546 800
rect 485686 0 485742 800
rect 486882 0 486938 800
rect 488078 0 488134 800
rect 489274 0 489330 800
rect 490470 0 490526 800
rect 491666 0 491722 800
rect 492862 0 492918 800
rect 494058 0 494114 800
rect 495254 0 495310 800
rect 496450 0 496506 800
rect 497646 0 497702 800
rect 498842 0 498898 800
rect 500038 0 500094 800
rect 501234 0 501290 800
rect 502430 0 502486 800
rect 503626 0 503682 800
rect 504822 0 504878 800
rect 506018 0 506074 800
rect 507214 0 507270 800
rect 508410 0 508466 800
rect 509606 0 509662 800
rect 510802 0 510858 800
rect 511998 0 512054 800
rect 513194 0 513250 800
rect 514390 0 514446 800
rect 515586 0 515642 800
rect 516782 0 516838 800
rect 517978 0 518034 800
rect 519174 0 519230 800
rect 520370 0 520426 800
rect 521566 0 521622 800
rect 522762 0 522818 800
rect 523958 0 524014 800
rect 525154 0 525210 800
rect 526350 0 526406 800
rect 527546 0 527602 800
rect 528742 0 528798 800
rect 529938 0 529994 800
rect 531134 0 531190 800
rect 532330 0 532386 800
rect 533526 0 533582 800
rect 534722 0 534778 800
rect 535918 0 535974 800
rect 537114 0 537170 800
rect 538310 0 538366 800
rect 539506 0 539562 800
rect 540702 0 540758 800
rect 541898 0 541954 800
rect 543094 0 543150 800
rect 544290 0 544346 800
rect 545486 0 545542 800
rect 546682 0 546738 800
rect 547878 0 547934 800
rect 549074 0 549130 800
rect 550270 0 550326 800
rect 551466 0 551522 800
rect 552662 0 552718 800
rect 553858 0 553914 800
<< obsm2 >>
rect 1582 499144 4838 499594
rect 5006 499144 9622 499594
rect 9790 499144 14406 499594
rect 14574 499144 19190 499594
rect 19358 499144 23974 499594
rect 24142 499144 28758 499594
rect 28926 499144 33542 499594
rect 33710 499144 38326 499594
rect 38494 499144 43110 499594
rect 43278 499144 47894 499594
rect 48062 499144 52678 499594
rect 52846 499144 57462 499594
rect 57630 499144 62246 499594
rect 62414 499144 67030 499594
rect 67198 499144 71814 499594
rect 71982 499144 76598 499594
rect 76766 499144 81382 499594
rect 81550 499144 86166 499594
rect 86334 499144 90950 499594
rect 91118 499144 95734 499594
rect 95902 499144 100518 499594
rect 100686 499144 105302 499594
rect 105470 499144 110086 499594
rect 110254 499144 114870 499594
rect 115038 499144 119654 499594
rect 119822 499144 124438 499594
rect 124606 499144 129222 499594
rect 129390 499144 134006 499594
rect 134174 499144 138790 499594
rect 138958 499144 143574 499594
rect 143742 499144 148358 499594
rect 148526 499144 153142 499594
rect 153310 499144 157926 499594
rect 158094 499144 162710 499594
rect 162878 499144 167494 499594
rect 167662 499144 172278 499594
rect 172446 499144 177062 499594
rect 177230 499144 181846 499594
rect 182014 499144 186630 499594
rect 186798 499144 191414 499594
rect 191582 499144 196198 499594
rect 196366 499144 200982 499594
rect 201150 499144 205766 499594
rect 205934 499144 210550 499594
rect 210718 499144 215334 499594
rect 215502 499144 220118 499594
rect 220286 499144 224902 499594
rect 225070 499144 229686 499594
rect 229854 499144 234470 499594
rect 234638 499144 239254 499594
rect 239422 499144 244038 499594
rect 244206 499144 248822 499594
rect 248990 499144 253606 499594
rect 253774 499144 258390 499594
rect 258558 499144 263174 499594
rect 263342 499144 267958 499594
rect 268126 499144 272742 499594
rect 272910 499144 277526 499594
rect 277694 499144 282310 499594
rect 282478 499144 287094 499594
rect 287262 499144 291878 499594
rect 292046 499144 296662 499594
rect 296830 499144 301446 499594
rect 301614 499144 306230 499594
rect 306398 499144 311014 499594
rect 311182 499144 315798 499594
rect 315966 499144 320582 499594
rect 320750 499144 325366 499594
rect 325534 499144 330150 499594
rect 330318 499144 334934 499594
rect 335102 499144 339718 499594
rect 339886 499144 344502 499594
rect 344670 499144 349286 499594
rect 349454 499144 354070 499594
rect 354238 499144 358854 499594
rect 359022 499144 363638 499594
rect 363806 499144 368422 499594
rect 368590 499144 373206 499594
rect 373374 499144 377990 499594
rect 378158 499144 382774 499594
rect 382942 499144 387558 499594
rect 387726 499144 392342 499594
rect 392510 499144 397126 499594
rect 397294 499144 401910 499594
rect 402078 499144 406694 499594
rect 406862 499144 411478 499594
rect 411646 499144 416262 499594
rect 416430 499144 421046 499594
rect 421214 499144 425830 499594
rect 425998 499144 430614 499594
rect 430782 499144 435398 499594
rect 435566 499144 440182 499594
rect 440350 499144 444966 499594
rect 445134 499144 449750 499594
rect 449918 499144 454534 499594
rect 454702 499144 459318 499594
rect 459486 499144 464102 499594
rect 464270 499144 468886 499594
rect 469054 499144 473670 499594
rect 473838 499144 478454 499594
rect 478622 499144 483238 499594
rect 483406 499144 488022 499594
rect 488190 499144 492806 499594
rect 492974 499144 497590 499594
rect 497758 499144 502374 499594
rect 502542 499144 507158 499594
rect 507326 499144 511942 499594
rect 512110 499144 516726 499594
rect 516894 499144 521510 499594
rect 521678 499144 526294 499594
rect 526462 499144 531078 499594
rect 531246 499144 535862 499594
rect 536030 499144 540646 499594
rect 540814 499144 545430 499594
rect 545598 499144 550214 499594
rect 550382 499144 554998 499594
rect 555166 499144 558512 499594
rect 1582 856 558512 499144
rect 1582 138 6034 856
rect 6202 138 7230 856
rect 7398 138 8426 856
rect 8594 138 9622 856
rect 9790 138 10818 856
rect 10986 138 12014 856
rect 12182 138 13210 856
rect 13378 138 14406 856
rect 14574 138 15602 856
rect 15770 138 16798 856
rect 16966 138 17994 856
rect 18162 138 19190 856
rect 19358 138 20386 856
rect 20554 138 21582 856
rect 21750 138 22778 856
rect 22946 138 23974 856
rect 24142 138 25170 856
rect 25338 138 26366 856
rect 26534 138 27562 856
rect 27730 138 28758 856
rect 28926 138 29954 856
rect 30122 138 31150 856
rect 31318 138 32346 856
rect 32514 138 33542 856
rect 33710 138 34738 856
rect 34906 138 35934 856
rect 36102 138 37130 856
rect 37298 138 38326 856
rect 38494 138 39522 856
rect 39690 138 40718 856
rect 40886 138 41914 856
rect 42082 138 43110 856
rect 43278 138 44306 856
rect 44474 138 45502 856
rect 45670 138 46698 856
rect 46866 138 47894 856
rect 48062 138 49090 856
rect 49258 138 50286 856
rect 50454 138 51482 856
rect 51650 138 52678 856
rect 52846 138 53874 856
rect 54042 138 55070 856
rect 55238 138 56266 856
rect 56434 138 57462 856
rect 57630 138 58658 856
rect 58826 138 59854 856
rect 60022 138 61050 856
rect 61218 138 62246 856
rect 62414 138 63442 856
rect 63610 138 64638 856
rect 64806 138 65834 856
rect 66002 138 67030 856
rect 67198 138 68226 856
rect 68394 138 69422 856
rect 69590 138 70618 856
rect 70786 138 71814 856
rect 71982 138 73010 856
rect 73178 138 74206 856
rect 74374 138 75402 856
rect 75570 138 76598 856
rect 76766 138 77794 856
rect 77962 138 78990 856
rect 79158 138 80186 856
rect 80354 138 81382 856
rect 81550 138 82578 856
rect 82746 138 83774 856
rect 83942 138 84970 856
rect 85138 138 86166 856
rect 86334 138 87362 856
rect 87530 138 88558 856
rect 88726 138 89754 856
rect 89922 138 90950 856
rect 91118 138 92146 856
rect 92314 138 93342 856
rect 93510 138 94538 856
rect 94706 138 95734 856
rect 95902 138 96930 856
rect 97098 138 98126 856
rect 98294 138 99322 856
rect 99490 138 100518 856
rect 100686 138 101714 856
rect 101882 138 102910 856
rect 103078 138 104106 856
rect 104274 138 105302 856
rect 105470 138 106498 856
rect 106666 138 107694 856
rect 107862 138 108890 856
rect 109058 138 110086 856
rect 110254 138 111282 856
rect 111450 138 112478 856
rect 112646 138 113674 856
rect 113842 138 114870 856
rect 115038 138 116066 856
rect 116234 138 117262 856
rect 117430 138 118458 856
rect 118626 138 119654 856
rect 119822 138 120850 856
rect 121018 138 122046 856
rect 122214 138 123242 856
rect 123410 138 124438 856
rect 124606 138 125634 856
rect 125802 138 126830 856
rect 126998 138 128026 856
rect 128194 138 129222 856
rect 129390 138 130418 856
rect 130586 138 131614 856
rect 131782 138 132810 856
rect 132978 138 134006 856
rect 134174 138 135202 856
rect 135370 138 136398 856
rect 136566 138 137594 856
rect 137762 138 138790 856
rect 138958 138 139986 856
rect 140154 138 141182 856
rect 141350 138 142378 856
rect 142546 138 143574 856
rect 143742 138 144770 856
rect 144938 138 145966 856
rect 146134 138 147162 856
rect 147330 138 148358 856
rect 148526 138 149554 856
rect 149722 138 150750 856
rect 150918 138 151946 856
rect 152114 138 153142 856
rect 153310 138 154338 856
rect 154506 138 155534 856
rect 155702 138 156730 856
rect 156898 138 157926 856
rect 158094 138 159122 856
rect 159290 138 160318 856
rect 160486 138 161514 856
rect 161682 138 162710 856
rect 162878 138 163906 856
rect 164074 138 165102 856
rect 165270 138 166298 856
rect 166466 138 167494 856
rect 167662 138 168690 856
rect 168858 138 169886 856
rect 170054 138 171082 856
rect 171250 138 172278 856
rect 172446 138 173474 856
rect 173642 138 174670 856
rect 174838 138 175866 856
rect 176034 138 177062 856
rect 177230 138 178258 856
rect 178426 138 179454 856
rect 179622 138 180650 856
rect 180818 138 181846 856
rect 182014 138 183042 856
rect 183210 138 184238 856
rect 184406 138 185434 856
rect 185602 138 186630 856
rect 186798 138 187826 856
rect 187994 138 189022 856
rect 189190 138 190218 856
rect 190386 138 191414 856
rect 191582 138 192610 856
rect 192778 138 193806 856
rect 193974 138 195002 856
rect 195170 138 196198 856
rect 196366 138 197394 856
rect 197562 138 198590 856
rect 198758 138 199786 856
rect 199954 138 200982 856
rect 201150 138 202178 856
rect 202346 138 203374 856
rect 203542 138 204570 856
rect 204738 138 205766 856
rect 205934 138 206962 856
rect 207130 138 208158 856
rect 208326 138 209354 856
rect 209522 138 210550 856
rect 210718 138 211746 856
rect 211914 138 212942 856
rect 213110 138 214138 856
rect 214306 138 215334 856
rect 215502 138 216530 856
rect 216698 138 217726 856
rect 217894 138 218922 856
rect 219090 138 220118 856
rect 220286 138 221314 856
rect 221482 138 222510 856
rect 222678 138 223706 856
rect 223874 138 224902 856
rect 225070 138 226098 856
rect 226266 138 227294 856
rect 227462 138 228490 856
rect 228658 138 229686 856
rect 229854 138 230882 856
rect 231050 138 232078 856
rect 232246 138 233274 856
rect 233442 138 234470 856
rect 234638 138 235666 856
rect 235834 138 236862 856
rect 237030 138 238058 856
rect 238226 138 239254 856
rect 239422 138 240450 856
rect 240618 138 241646 856
rect 241814 138 242842 856
rect 243010 138 244038 856
rect 244206 138 245234 856
rect 245402 138 246430 856
rect 246598 138 247626 856
rect 247794 138 248822 856
rect 248990 138 250018 856
rect 250186 138 251214 856
rect 251382 138 252410 856
rect 252578 138 253606 856
rect 253774 138 254802 856
rect 254970 138 255998 856
rect 256166 138 257194 856
rect 257362 138 258390 856
rect 258558 138 259586 856
rect 259754 138 260782 856
rect 260950 138 261978 856
rect 262146 138 263174 856
rect 263342 138 264370 856
rect 264538 138 265566 856
rect 265734 138 266762 856
rect 266930 138 267958 856
rect 268126 138 269154 856
rect 269322 138 270350 856
rect 270518 138 271546 856
rect 271714 138 272742 856
rect 272910 138 273938 856
rect 274106 138 275134 856
rect 275302 138 276330 856
rect 276498 138 277526 856
rect 277694 138 278722 856
rect 278890 138 279918 856
rect 280086 138 281114 856
rect 281282 138 282310 856
rect 282478 138 283506 856
rect 283674 138 284702 856
rect 284870 138 285898 856
rect 286066 138 287094 856
rect 287262 138 288290 856
rect 288458 138 289486 856
rect 289654 138 290682 856
rect 290850 138 291878 856
rect 292046 138 293074 856
rect 293242 138 294270 856
rect 294438 138 295466 856
rect 295634 138 296662 856
rect 296830 138 297858 856
rect 298026 138 299054 856
rect 299222 138 300250 856
rect 300418 138 301446 856
rect 301614 138 302642 856
rect 302810 138 303838 856
rect 304006 138 305034 856
rect 305202 138 306230 856
rect 306398 138 307426 856
rect 307594 138 308622 856
rect 308790 138 309818 856
rect 309986 138 311014 856
rect 311182 138 312210 856
rect 312378 138 313406 856
rect 313574 138 314602 856
rect 314770 138 315798 856
rect 315966 138 316994 856
rect 317162 138 318190 856
rect 318358 138 319386 856
rect 319554 138 320582 856
rect 320750 138 321778 856
rect 321946 138 322974 856
rect 323142 138 324170 856
rect 324338 138 325366 856
rect 325534 138 326562 856
rect 326730 138 327758 856
rect 327926 138 328954 856
rect 329122 138 330150 856
rect 330318 138 331346 856
rect 331514 138 332542 856
rect 332710 138 333738 856
rect 333906 138 334934 856
rect 335102 138 336130 856
rect 336298 138 337326 856
rect 337494 138 338522 856
rect 338690 138 339718 856
rect 339886 138 340914 856
rect 341082 138 342110 856
rect 342278 138 343306 856
rect 343474 138 344502 856
rect 344670 138 345698 856
rect 345866 138 346894 856
rect 347062 138 348090 856
rect 348258 138 349286 856
rect 349454 138 350482 856
rect 350650 138 351678 856
rect 351846 138 352874 856
rect 353042 138 354070 856
rect 354238 138 355266 856
rect 355434 138 356462 856
rect 356630 138 357658 856
rect 357826 138 358854 856
rect 359022 138 360050 856
rect 360218 138 361246 856
rect 361414 138 362442 856
rect 362610 138 363638 856
rect 363806 138 364834 856
rect 365002 138 366030 856
rect 366198 138 367226 856
rect 367394 138 368422 856
rect 368590 138 369618 856
rect 369786 138 370814 856
rect 370982 138 372010 856
rect 372178 138 373206 856
rect 373374 138 374402 856
rect 374570 138 375598 856
rect 375766 138 376794 856
rect 376962 138 377990 856
rect 378158 138 379186 856
rect 379354 138 380382 856
rect 380550 138 381578 856
rect 381746 138 382774 856
rect 382942 138 383970 856
rect 384138 138 385166 856
rect 385334 138 386362 856
rect 386530 138 387558 856
rect 387726 138 388754 856
rect 388922 138 389950 856
rect 390118 138 391146 856
rect 391314 138 392342 856
rect 392510 138 393538 856
rect 393706 138 394734 856
rect 394902 138 395930 856
rect 396098 138 397126 856
rect 397294 138 398322 856
rect 398490 138 399518 856
rect 399686 138 400714 856
rect 400882 138 401910 856
rect 402078 138 403106 856
rect 403274 138 404302 856
rect 404470 138 405498 856
rect 405666 138 406694 856
rect 406862 138 407890 856
rect 408058 138 409086 856
rect 409254 138 410282 856
rect 410450 138 411478 856
rect 411646 138 412674 856
rect 412842 138 413870 856
rect 414038 138 415066 856
rect 415234 138 416262 856
rect 416430 138 417458 856
rect 417626 138 418654 856
rect 418822 138 419850 856
rect 420018 138 421046 856
rect 421214 138 422242 856
rect 422410 138 423438 856
rect 423606 138 424634 856
rect 424802 138 425830 856
rect 425998 138 427026 856
rect 427194 138 428222 856
rect 428390 138 429418 856
rect 429586 138 430614 856
rect 430782 138 431810 856
rect 431978 138 433006 856
rect 433174 138 434202 856
rect 434370 138 435398 856
rect 435566 138 436594 856
rect 436762 138 437790 856
rect 437958 138 438986 856
rect 439154 138 440182 856
rect 440350 138 441378 856
rect 441546 138 442574 856
rect 442742 138 443770 856
rect 443938 138 444966 856
rect 445134 138 446162 856
rect 446330 138 447358 856
rect 447526 138 448554 856
rect 448722 138 449750 856
rect 449918 138 450946 856
rect 451114 138 452142 856
rect 452310 138 453338 856
rect 453506 138 454534 856
rect 454702 138 455730 856
rect 455898 138 456926 856
rect 457094 138 458122 856
rect 458290 138 459318 856
rect 459486 138 460514 856
rect 460682 138 461710 856
rect 461878 138 462906 856
rect 463074 138 464102 856
rect 464270 138 465298 856
rect 465466 138 466494 856
rect 466662 138 467690 856
rect 467858 138 468886 856
rect 469054 138 470082 856
rect 470250 138 471278 856
rect 471446 138 472474 856
rect 472642 138 473670 856
rect 473838 138 474866 856
rect 475034 138 476062 856
rect 476230 138 477258 856
rect 477426 138 478454 856
rect 478622 138 479650 856
rect 479818 138 480846 856
rect 481014 138 482042 856
rect 482210 138 483238 856
rect 483406 138 484434 856
rect 484602 138 485630 856
rect 485798 138 486826 856
rect 486994 138 488022 856
rect 488190 138 489218 856
rect 489386 138 490414 856
rect 490582 138 491610 856
rect 491778 138 492806 856
rect 492974 138 494002 856
rect 494170 138 495198 856
rect 495366 138 496394 856
rect 496562 138 497590 856
rect 497758 138 498786 856
rect 498954 138 499982 856
rect 500150 138 501178 856
rect 501346 138 502374 856
rect 502542 138 503570 856
rect 503738 138 504766 856
rect 504934 138 505962 856
rect 506130 138 507158 856
rect 507326 138 508354 856
rect 508522 138 509550 856
rect 509718 138 510746 856
rect 510914 138 511942 856
rect 512110 138 513138 856
rect 513306 138 514334 856
rect 514502 138 515530 856
rect 515698 138 516726 856
rect 516894 138 517922 856
rect 518090 138 519118 856
rect 519286 138 520314 856
rect 520482 138 521510 856
rect 521678 138 522706 856
rect 522874 138 523902 856
rect 524070 138 525098 856
rect 525266 138 526294 856
rect 526462 138 527490 856
rect 527658 138 528686 856
rect 528854 138 529882 856
rect 530050 138 531078 856
rect 531246 138 532274 856
rect 532442 138 533470 856
rect 533638 138 534666 856
rect 534834 138 535862 856
rect 536030 138 537058 856
rect 537226 138 538254 856
rect 538422 138 539450 856
rect 539618 138 540646 856
rect 540814 138 541842 856
rect 542010 138 543038 856
rect 543206 138 544234 856
rect 544402 138 545430 856
rect 545598 138 546626 856
rect 546794 138 547822 856
rect 547990 138 549018 856
rect 549186 138 550214 856
rect 550382 138 551410 856
rect 551578 138 552606 856
rect 552774 138 553802 856
rect 553970 138 558512 856
<< metal3 >>
rect 0 494912 800 495032
rect 559200 493824 560000 493944
rect 0 485664 800 485784
rect 559200 484440 560000 484560
rect 0 476416 800 476536
rect 559200 475056 560000 475176
rect 0 467168 800 467288
rect 559200 465672 560000 465792
rect 0 457920 800 458040
rect 559200 456288 560000 456408
rect 0 448672 800 448792
rect 559200 446904 560000 447024
rect 0 439424 800 439544
rect 559200 437520 560000 437640
rect 0 430176 800 430296
rect 559200 428136 560000 428256
rect 0 420928 800 421048
rect 559200 418752 560000 418872
rect 0 411680 800 411800
rect 559200 409368 560000 409488
rect 0 402432 800 402552
rect 559200 399984 560000 400104
rect 0 393184 800 393304
rect 559200 390600 560000 390720
rect 0 383936 800 384056
rect 559200 381216 560000 381336
rect 0 374688 800 374808
rect 559200 371832 560000 371952
rect 0 365440 800 365560
rect 559200 362448 560000 362568
rect 0 356192 800 356312
rect 559200 353064 560000 353184
rect 0 346944 800 347064
rect 559200 343680 560000 343800
rect 0 337696 800 337816
rect 559200 334296 560000 334416
rect 0 328448 800 328568
rect 559200 324912 560000 325032
rect 0 319200 800 319320
rect 559200 315528 560000 315648
rect 0 309952 800 310072
rect 559200 306144 560000 306264
rect 0 300704 800 300824
rect 559200 296760 560000 296880
rect 0 291456 800 291576
rect 559200 287376 560000 287496
rect 0 282208 800 282328
rect 559200 277992 560000 278112
rect 0 272960 800 273080
rect 559200 268608 560000 268728
rect 0 263712 800 263832
rect 559200 259224 560000 259344
rect 0 254464 800 254584
rect 559200 249840 560000 249960
rect 0 245216 800 245336
rect 559200 240456 560000 240576
rect 0 235968 800 236088
rect 559200 231072 560000 231192
rect 0 226720 800 226840
rect 559200 221688 560000 221808
rect 0 217472 800 217592
rect 559200 212304 560000 212424
rect 0 208224 800 208344
rect 559200 202920 560000 203040
rect 0 198976 800 199096
rect 559200 193536 560000 193656
rect 0 189728 800 189848
rect 559200 184152 560000 184272
rect 0 180480 800 180600
rect 559200 174768 560000 174888
rect 0 171232 800 171352
rect 559200 165384 560000 165504
rect 0 161984 800 162104
rect 559200 156000 560000 156120
rect 0 152736 800 152856
rect 559200 146616 560000 146736
rect 0 143488 800 143608
rect 559200 137232 560000 137352
rect 0 134240 800 134360
rect 559200 127848 560000 127968
rect 0 124992 800 125112
rect 559200 118464 560000 118584
rect 0 115744 800 115864
rect 559200 109080 560000 109200
rect 0 106496 800 106616
rect 559200 99696 560000 99816
rect 0 97248 800 97368
rect 559200 90312 560000 90432
rect 0 88000 800 88120
rect 559200 80928 560000 81048
rect 0 78752 800 78872
rect 559200 71544 560000 71664
rect 0 69504 800 69624
rect 559200 62160 560000 62280
rect 0 60256 800 60376
rect 559200 52776 560000 52896
rect 0 51008 800 51128
rect 559200 43392 560000 43512
rect 0 41760 800 41880
rect 559200 34008 560000 34128
rect 0 32512 800 32632
rect 559200 24624 560000 24744
rect 0 23264 800 23384
rect 559200 15240 560000 15360
rect 0 14016 800 14136
rect 559200 5856 560000 5976
rect 0 4768 800 4888
<< obsm3 >>
rect 800 495112 559200 499085
rect 880 494832 559200 495112
rect 800 494024 559200 494832
rect 800 493744 559120 494024
rect 800 485864 559200 493744
rect 880 485584 559200 485864
rect 800 484640 559200 485584
rect 800 484360 559120 484640
rect 800 476616 559200 484360
rect 880 476336 559200 476616
rect 800 475256 559200 476336
rect 800 474976 559120 475256
rect 800 467368 559200 474976
rect 880 467088 559200 467368
rect 800 465872 559200 467088
rect 800 465592 559120 465872
rect 800 458120 559200 465592
rect 880 457840 559200 458120
rect 800 456488 559200 457840
rect 800 456208 559120 456488
rect 800 448872 559200 456208
rect 880 448592 559200 448872
rect 800 447104 559200 448592
rect 800 446824 559120 447104
rect 800 439624 559200 446824
rect 880 439344 559200 439624
rect 800 437720 559200 439344
rect 800 437440 559120 437720
rect 800 430376 559200 437440
rect 880 430096 559200 430376
rect 800 428336 559200 430096
rect 800 428056 559120 428336
rect 800 421128 559200 428056
rect 880 420848 559200 421128
rect 800 418952 559200 420848
rect 800 418672 559120 418952
rect 800 411880 559200 418672
rect 880 411600 559200 411880
rect 800 409568 559200 411600
rect 800 409288 559120 409568
rect 800 402632 559200 409288
rect 880 402352 559200 402632
rect 800 400184 559200 402352
rect 800 399904 559120 400184
rect 800 393384 559200 399904
rect 880 393104 559200 393384
rect 800 390800 559200 393104
rect 800 390520 559120 390800
rect 800 384136 559200 390520
rect 880 383856 559200 384136
rect 800 381416 559200 383856
rect 800 381136 559120 381416
rect 800 374888 559200 381136
rect 880 374608 559200 374888
rect 800 372032 559200 374608
rect 800 371752 559120 372032
rect 800 365640 559200 371752
rect 880 365360 559200 365640
rect 800 362648 559200 365360
rect 800 362368 559120 362648
rect 800 356392 559200 362368
rect 880 356112 559200 356392
rect 800 353264 559200 356112
rect 800 352984 559120 353264
rect 800 347144 559200 352984
rect 880 346864 559200 347144
rect 800 343880 559200 346864
rect 800 343600 559120 343880
rect 800 337896 559200 343600
rect 880 337616 559200 337896
rect 800 334496 559200 337616
rect 800 334216 559120 334496
rect 800 328648 559200 334216
rect 880 328368 559200 328648
rect 800 325112 559200 328368
rect 800 324832 559120 325112
rect 800 319400 559200 324832
rect 880 319120 559200 319400
rect 800 315728 559200 319120
rect 800 315448 559120 315728
rect 800 310152 559200 315448
rect 880 309872 559200 310152
rect 800 306344 559200 309872
rect 800 306064 559120 306344
rect 800 300904 559200 306064
rect 880 300624 559200 300904
rect 800 296960 559200 300624
rect 800 296680 559120 296960
rect 800 291656 559200 296680
rect 880 291376 559200 291656
rect 800 287576 559200 291376
rect 800 287296 559120 287576
rect 800 282408 559200 287296
rect 880 282128 559200 282408
rect 800 278192 559200 282128
rect 800 277912 559120 278192
rect 800 273160 559200 277912
rect 880 272880 559200 273160
rect 800 268808 559200 272880
rect 800 268528 559120 268808
rect 800 263912 559200 268528
rect 880 263632 559200 263912
rect 800 259424 559200 263632
rect 800 259144 559120 259424
rect 800 254664 559200 259144
rect 880 254384 559200 254664
rect 800 250040 559200 254384
rect 800 249760 559120 250040
rect 800 245416 559200 249760
rect 880 245136 559200 245416
rect 800 240656 559200 245136
rect 800 240376 559120 240656
rect 800 236168 559200 240376
rect 880 235888 559200 236168
rect 800 231272 559200 235888
rect 800 230992 559120 231272
rect 800 226920 559200 230992
rect 880 226640 559200 226920
rect 800 221888 559200 226640
rect 800 221608 559120 221888
rect 800 217672 559200 221608
rect 880 217392 559200 217672
rect 800 212504 559200 217392
rect 800 212224 559120 212504
rect 800 208424 559200 212224
rect 880 208144 559200 208424
rect 800 203120 559200 208144
rect 800 202840 559120 203120
rect 800 199176 559200 202840
rect 880 198896 559200 199176
rect 800 193736 559200 198896
rect 800 193456 559120 193736
rect 800 189928 559200 193456
rect 880 189648 559200 189928
rect 800 184352 559200 189648
rect 800 184072 559120 184352
rect 800 180680 559200 184072
rect 880 180400 559200 180680
rect 800 174968 559200 180400
rect 800 174688 559120 174968
rect 800 171432 559200 174688
rect 880 171152 559200 171432
rect 800 165584 559200 171152
rect 800 165304 559120 165584
rect 800 162184 559200 165304
rect 880 161904 559200 162184
rect 800 156200 559200 161904
rect 800 155920 559120 156200
rect 800 152936 559200 155920
rect 880 152656 559200 152936
rect 800 146816 559200 152656
rect 800 146536 559120 146816
rect 800 143688 559200 146536
rect 880 143408 559200 143688
rect 800 137432 559200 143408
rect 800 137152 559120 137432
rect 800 134440 559200 137152
rect 880 134160 559200 134440
rect 800 128048 559200 134160
rect 800 127768 559120 128048
rect 800 125192 559200 127768
rect 880 124912 559200 125192
rect 800 118664 559200 124912
rect 800 118384 559120 118664
rect 800 115944 559200 118384
rect 880 115664 559200 115944
rect 800 109280 559200 115664
rect 800 109000 559120 109280
rect 800 106696 559200 109000
rect 880 106416 559200 106696
rect 800 99896 559200 106416
rect 800 99616 559120 99896
rect 800 97448 559200 99616
rect 880 97168 559200 97448
rect 800 90512 559200 97168
rect 800 90232 559120 90512
rect 800 88200 559200 90232
rect 880 87920 559200 88200
rect 800 81128 559200 87920
rect 800 80848 559120 81128
rect 800 78952 559200 80848
rect 880 78672 559200 78952
rect 800 71744 559200 78672
rect 800 71464 559120 71744
rect 800 69704 559200 71464
rect 880 69424 559200 69704
rect 800 62360 559200 69424
rect 800 62080 559120 62360
rect 800 60456 559200 62080
rect 880 60176 559200 60456
rect 800 52976 559200 60176
rect 800 52696 559120 52976
rect 800 51208 559200 52696
rect 880 50928 559200 51208
rect 800 43592 559200 50928
rect 800 43312 559120 43592
rect 800 41960 559200 43312
rect 880 41680 559200 41960
rect 800 34208 559200 41680
rect 800 33928 559120 34208
rect 800 32712 559200 33928
rect 880 32432 559200 32712
rect 800 24824 559200 32432
rect 800 24544 559120 24824
rect 800 23464 559200 24544
rect 880 23184 559200 23464
rect 800 15440 559200 23184
rect 800 15160 559120 15440
rect 800 14216 559200 15160
rect 880 13936 559200 14216
rect 800 6056 559200 13936
rect 800 5776 559120 6056
rect 800 4968 559200 5776
rect 880 4688 559200 4968
rect 800 443 559200 4688
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
rect 34928 2128 35248 497808
rect 50288 2128 50608 497808
rect 65648 2128 65968 497808
rect 81008 2128 81328 497808
rect 96368 2128 96688 497808
rect 111728 2128 112048 497808
rect 127088 2128 127408 497808
rect 142448 2128 142768 497808
rect 157808 2128 158128 497808
rect 173168 2128 173488 497808
rect 188528 2128 188848 497808
rect 203888 2128 204208 497808
rect 219248 2128 219568 497808
rect 234608 2128 234928 497808
rect 249968 2128 250288 497808
rect 265328 2128 265648 497808
rect 280688 2128 281008 497808
rect 296048 2128 296368 497808
rect 311408 2128 311728 497808
rect 326768 2128 327088 497808
rect 342128 2128 342448 497808
rect 357488 2128 357808 497808
rect 372848 2128 373168 497808
rect 388208 2128 388528 497808
rect 403568 2128 403888 497808
rect 418928 2128 419248 497808
rect 434288 2128 434608 497808
rect 449648 2128 449968 497808
rect 465008 2128 465328 497808
rect 480368 2128 480688 497808
rect 495728 2128 496048 497808
rect 511088 2128 511408 497808
rect 526448 2128 526768 497808
rect 541808 2128 542128 497808
rect 557168 2128 557488 497808
<< obsm4 >>
rect 17539 497888 546237 499085
rect 17539 2048 19488 497888
rect 19968 2048 34848 497888
rect 35328 2048 50208 497888
rect 50688 2048 65568 497888
rect 66048 2048 80928 497888
rect 81408 2048 96288 497888
rect 96768 2048 111648 497888
rect 112128 2048 127008 497888
rect 127488 2048 142368 497888
rect 142848 2048 157728 497888
rect 158208 2048 173088 497888
rect 173568 2048 188448 497888
rect 188928 2048 203808 497888
rect 204288 2048 219168 497888
rect 219648 2048 234528 497888
rect 235008 2048 249888 497888
rect 250368 2048 265248 497888
rect 265728 2048 280608 497888
rect 281088 2048 295968 497888
rect 296448 2048 311328 497888
rect 311808 2048 326688 497888
rect 327168 2048 342048 497888
rect 342528 2048 357408 497888
rect 357888 2048 372768 497888
rect 373248 2048 388128 497888
rect 388608 2048 403488 497888
rect 403968 2048 418848 497888
rect 419328 2048 434208 497888
rect 434688 2048 449568 497888
rect 450048 2048 464928 497888
rect 465408 2048 480288 497888
rect 480768 2048 495648 497888
rect 496128 2048 511008 497888
rect 511488 2048 526368 497888
rect 526848 2048 541728 497888
rect 542208 2048 546237 497888
rect 17539 579 546237 2048
<< labels >>
rlabel metal3 s 559200 428136 560000 428256 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 397182 499200 397238 500000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 401966 499200 402022 500000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 406750 499200 406806 500000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 411534 499200 411590 500000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 416318 499200 416374 500000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 421102 499200 421158 500000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 425886 499200 425942 500000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 393184 800 393304 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 402432 800 402552 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 411680 800 411800 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 559200 437520 560000 437640 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 420928 800 421048 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 430176 800 430296 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 439424 800 439544 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 448672 800 448792 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 457920 800 458040 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 467168 800 467288 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 476416 800 476536 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 485664 800 485784 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 494912 800 495032 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 559200 446904 560000 447024 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 559200 456288 560000 456408 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 559200 465672 560000 465792 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 559200 475056 560000 475176 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 559200 484440 560000 484560 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 559200 493824 560000 493944 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 387614 499200 387670 500000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 392398 499200 392454 500000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 290738 0 290794 800 6 instrMgmt_addr[0]
port 30 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 instrMgmt_addr[1]
port 31 nsew signal output
rlabel metal2 s 293130 0 293186 800 6 instrMgmt_addr[2]
port 32 nsew signal output
rlabel metal2 s 294326 0 294382 800 6 instrMgmt_addr[3]
port 33 nsew signal output
rlabel metal2 s 295522 0 295578 800 6 instrMgmt_addr[4]
port 34 nsew signal output
rlabel metal2 s 296718 0 296774 800 6 instrMgmt_addr[5]
port 35 nsew signal output
rlabel metal2 s 297914 0 297970 800 6 instrMgmt_addr[6]
port 36 nsew signal output
rlabel metal2 s 299110 0 299166 800 6 instrMgmt_addr[7]
port 37 nsew signal output
rlabel metal2 s 300306 0 300362 800 6 instrMgmt_addr[8]
port 38 nsew signal output
rlabel metal2 s 454590 0 454646 800 6 instrMgmt_ce
port 39 nsew signal output
rlabel metal2 s 301502 0 301558 800 6 instrMgmt_dataIn[0]
port 40 nsew signal input
rlabel metal2 s 313462 0 313518 800 6 instrMgmt_dataIn[10]
port 41 nsew signal input
rlabel metal2 s 314658 0 314714 800 6 instrMgmt_dataIn[11]
port 42 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 instrMgmt_dataIn[12]
port 43 nsew signal input
rlabel metal2 s 317050 0 317106 800 6 instrMgmt_dataIn[13]
port 44 nsew signal input
rlabel metal2 s 318246 0 318302 800 6 instrMgmt_dataIn[14]
port 45 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 instrMgmt_dataIn[15]
port 46 nsew signal input
rlabel metal2 s 320638 0 320694 800 6 instrMgmt_dataIn[16]
port 47 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 instrMgmt_dataIn[17]
port 48 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 instrMgmt_dataIn[18]
port 49 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 instrMgmt_dataIn[19]
port 50 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 instrMgmt_dataIn[1]
port 51 nsew signal input
rlabel metal2 s 325422 0 325478 800 6 instrMgmt_dataIn[20]
port 52 nsew signal input
rlabel metal2 s 326618 0 326674 800 6 instrMgmt_dataIn[21]
port 53 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 instrMgmt_dataIn[22]
port 54 nsew signal input
rlabel metal2 s 329010 0 329066 800 6 instrMgmt_dataIn[23]
port 55 nsew signal input
rlabel metal2 s 330206 0 330262 800 6 instrMgmt_dataIn[24]
port 56 nsew signal input
rlabel metal2 s 331402 0 331458 800 6 instrMgmt_dataIn[25]
port 57 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 instrMgmt_dataIn[26]
port 58 nsew signal input
rlabel metal2 s 333794 0 333850 800 6 instrMgmt_dataIn[27]
port 59 nsew signal input
rlabel metal2 s 334990 0 335046 800 6 instrMgmt_dataIn[28]
port 60 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 instrMgmt_dataIn[29]
port 61 nsew signal input
rlabel metal2 s 303894 0 303950 800 6 instrMgmt_dataIn[2]
port 62 nsew signal input
rlabel metal2 s 337382 0 337438 800 6 instrMgmt_dataIn[30]
port 63 nsew signal input
rlabel metal2 s 338578 0 338634 800 6 instrMgmt_dataIn[31]
port 64 nsew signal input
rlabel metal2 s 339774 0 339830 800 6 instrMgmt_dataIn[32]
port 65 nsew signal input
rlabel metal2 s 340970 0 341026 800 6 instrMgmt_dataIn[33]
port 66 nsew signal input
rlabel metal2 s 342166 0 342222 800 6 instrMgmt_dataIn[34]
port 67 nsew signal input
rlabel metal2 s 343362 0 343418 800 6 instrMgmt_dataIn[35]
port 68 nsew signal input
rlabel metal2 s 344558 0 344614 800 6 instrMgmt_dataIn[36]
port 69 nsew signal input
rlabel metal2 s 345754 0 345810 800 6 instrMgmt_dataIn[37]
port 70 nsew signal input
rlabel metal2 s 346950 0 347006 800 6 instrMgmt_dataIn[38]
port 71 nsew signal input
rlabel metal2 s 348146 0 348202 800 6 instrMgmt_dataIn[39]
port 72 nsew signal input
rlabel metal2 s 305090 0 305146 800 6 instrMgmt_dataIn[3]
port 73 nsew signal input
rlabel metal2 s 349342 0 349398 800 6 instrMgmt_dataIn[40]
port 74 nsew signal input
rlabel metal2 s 350538 0 350594 800 6 instrMgmt_dataIn[41]
port 75 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 instrMgmt_dataIn[42]
port 76 nsew signal input
rlabel metal2 s 352930 0 352986 800 6 instrMgmt_dataIn[43]
port 77 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 instrMgmt_dataIn[44]
port 78 nsew signal input
rlabel metal2 s 355322 0 355378 800 6 instrMgmt_dataIn[45]
port 79 nsew signal input
rlabel metal2 s 356518 0 356574 800 6 instrMgmt_dataIn[46]
port 80 nsew signal input
rlabel metal2 s 357714 0 357770 800 6 instrMgmt_dataIn[47]
port 81 nsew signal input
rlabel metal2 s 358910 0 358966 800 6 instrMgmt_dataIn[48]
port 82 nsew signal input
rlabel metal2 s 360106 0 360162 800 6 instrMgmt_dataIn[49]
port 83 nsew signal input
rlabel metal2 s 306286 0 306342 800 6 instrMgmt_dataIn[4]
port 84 nsew signal input
rlabel metal2 s 361302 0 361358 800 6 instrMgmt_dataIn[50]
port 85 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 instrMgmt_dataIn[51]
port 86 nsew signal input
rlabel metal2 s 363694 0 363750 800 6 instrMgmt_dataIn[52]
port 87 nsew signal input
rlabel metal2 s 364890 0 364946 800 6 instrMgmt_dataIn[53]
port 88 nsew signal input
rlabel metal2 s 366086 0 366142 800 6 instrMgmt_dataIn[54]
port 89 nsew signal input
rlabel metal2 s 367282 0 367338 800 6 instrMgmt_dataIn[55]
port 90 nsew signal input
rlabel metal2 s 368478 0 368534 800 6 instrMgmt_dataIn[56]
port 91 nsew signal input
rlabel metal2 s 369674 0 369730 800 6 instrMgmt_dataIn[57]
port 92 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 instrMgmt_dataIn[58]
port 93 nsew signal input
rlabel metal2 s 372066 0 372122 800 6 instrMgmt_dataIn[59]
port 94 nsew signal input
rlabel metal2 s 307482 0 307538 800 6 instrMgmt_dataIn[5]
port 95 nsew signal input
rlabel metal2 s 373262 0 373318 800 6 instrMgmt_dataIn[60]
port 96 nsew signal input
rlabel metal2 s 374458 0 374514 800 6 instrMgmt_dataIn[61]
port 97 nsew signal input
rlabel metal2 s 375654 0 375710 800 6 instrMgmt_dataIn[62]
port 98 nsew signal input
rlabel metal2 s 376850 0 376906 800 6 instrMgmt_dataIn[63]
port 99 nsew signal input
rlabel metal2 s 308678 0 308734 800 6 instrMgmt_dataIn[6]
port 100 nsew signal input
rlabel metal2 s 309874 0 309930 800 6 instrMgmt_dataIn[7]
port 101 nsew signal input
rlabel metal2 s 311070 0 311126 800 6 instrMgmt_dataIn[8]
port 102 nsew signal input
rlabel metal2 s 312266 0 312322 800 6 instrMgmt_dataIn[9]
port 103 nsew signal input
rlabel metal2 s 378046 0 378102 800 6 instrMgmt_dataOut[0]
port 104 nsew signal output
rlabel metal2 s 390006 0 390062 800 6 instrMgmt_dataOut[10]
port 105 nsew signal output
rlabel metal2 s 391202 0 391258 800 6 instrMgmt_dataOut[11]
port 106 nsew signal output
rlabel metal2 s 392398 0 392454 800 6 instrMgmt_dataOut[12]
port 107 nsew signal output
rlabel metal2 s 393594 0 393650 800 6 instrMgmt_dataOut[13]
port 108 nsew signal output
rlabel metal2 s 394790 0 394846 800 6 instrMgmt_dataOut[14]
port 109 nsew signal output
rlabel metal2 s 395986 0 396042 800 6 instrMgmt_dataOut[15]
port 110 nsew signal output
rlabel metal2 s 397182 0 397238 800 6 instrMgmt_dataOut[16]
port 111 nsew signal output
rlabel metal2 s 398378 0 398434 800 6 instrMgmt_dataOut[17]
port 112 nsew signal output
rlabel metal2 s 399574 0 399630 800 6 instrMgmt_dataOut[18]
port 113 nsew signal output
rlabel metal2 s 400770 0 400826 800 6 instrMgmt_dataOut[19]
port 114 nsew signal output
rlabel metal2 s 379242 0 379298 800 6 instrMgmt_dataOut[1]
port 115 nsew signal output
rlabel metal2 s 401966 0 402022 800 6 instrMgmt_dataOut[20]
port 116 nsew signal output
rlabel metal2 s 403162 0 403218 800 6 instrMgmt_dataOut[21]
port 117 nsew signal output
rlabel metal2 s 404358 0 404414 800 6 instrMgmt_dataOut[22]
port 118 nsew signal output
rlabel metal2 s 405554 0 405610 800 6 instrMgmt_dataOut[23]
port 119 nsew signal output
rlabel metal2 s 406750 0 406806 800 6 instrMgmt_dataOut[24]
port 120 nsew signal output
rlabel metal2 s 407946 0 408002 800 6 instrMgmt_dataOut[25]
port 121 nsew signal output
rlabel metal2 s 409142 0 409198 800 6 instrMgmt_dataOut[26]
port 122 nsew signal output
rlabel metal2 s 410338 0 410394 800 6 instrMgmt_dataOut[27]
port 123 nsew signal output
rlabel metal2 s 411534 0 411590 800 6 instrMgmt_dataOut[28]
port 124 nsew signal output
rlabel metal2 s 412730 0 412786 800 6 instrMgmt_dataOut[29]
port 125 nsew signal output
rlabel metal2 s 380438 0 380494 800 6 instrMgmt_dataOut[2]
port 126 nsew signal output
rlabel metal2 s 413926 0 413982 800 6 instrMgmt_dataOut[30]
port 127 nsew signal output
rlabel metal2 s 415122 0 415178 800 6 instrMgmt_dataOut[31]
port 128 nsew signal output
rlabel metal2 s 416318 0 416374 800 6 instrMgmt_dataOut[32]
port 129 nsew signal output
rlabel metal2 s 417514 0 417570 800 6 instrMgmt_dataOut[33]
port 130 nsew signal output
rlabel metal2 s 418710 0 418766 800 6 instrMgmt_dataOut[34]
port 131 nsew signal output
rlabel metal2 s 419906 0 419962 800 6 instrMgmt_dataOut[35]
port 132 nsew signal output
rlabel metal2 s 421102 0 421158 800 6 instrMgmt_dataOut[36]
port 133 nsew signal output
rlabel metal2 s 422298 0 422354 800 6 instrMgmt_dataOut[37]
port 134 nsew signal output
rlabel metal2 s 423494 0 423550 800 6 instrMgmt_dataOut[38]
port 135 nsew signal output
rlabel metal2 s 424690 0 424746 800 6 instrMgmt_dataOut[39]
port 136 nsew signal output
rlabel metal2 s 381634 0 381690 800 6 instrMgmt_dataOut[3]
port 137 nsew signal output
rlabel metal2 s 425886 0 425942 800 6 instrMgmt_dataOut[40]
port 138 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 instrMgmt_dataOut[41]
port 139 nsew signal output
rlabel metal2 s 428278 0 428334 800 6 instrMgmt_dataOut[42]
port 140 nsew signal output
rlabel metal2 s 429474 0 429530 800 6 instrMgmt_dataOut[43]
port 141 nsew signal output
rlabel metal2 s 430670 0 430726 800 6 instrMgmt_dataOut[44]
port 142 nsew signal output
rlabel metal2 s 431866 0 431922 800 6 instrMgmt_dataOut[45]
port 143 nsew signal output
rlabel metal2 s 433062 0 433118 800 6 instrMgmt_dataOut[46]
port 144 nsew signal output
rlabel metal2 s 434258 0 434314 800 6 instrMgmt_dataOut[47]
port 145 nsew signal output
rlabel metal2 s 435454 0 435510 800 6 instrMgmt_dataOut[48]
port 146 nsew signal output
rlabel metal2 s 436650 0 436706 800 6 instrMgmt_dataOut[49]
port 147 nsew signal output
rlabel metal2 s 382830 0 382886 800 6 instrMgmt_dataOut[4]
port 148 nsew signal output
rlabel metal2 s 437846 0 437902 800 6 instrMgmt_dataOut[50]
port 149 nsew signal output
rlabel metal2 s 439042 0 439098 800 6 instrMgmt_dataOut[51]
port 150 nsew signal output
rlabel metal2 s 440238 0 440294 800 6 instrMgmt_dataOut[52]
port 151 nsew signal output
rlabel metal2 s 441434 0 441490 800 6 instrMgmt_dataOut[53]
port 152 nsew signal output
rlabel metal2 s 442630 0 442686 800 6 instrMgmt_dataOut[54]
port 153 nsew signal output
rlabel metal2 s 443826 0 443882 800 6 instrMgmt_dataOut[55]
port 154 nsew signal output
rlabel metal2 s 445022 0 445078 800 6 instrMgmt_dataOut[56]
port 155 nsew signal output
rlabel metal2 s 446218 0 446274 800 6 instrMgmt_dataOut[57]
port 156 nsew signal output
rlabel metal2 s 447414 0 447470 800 6 instrMgmt_dataOut[58]
port 157 nsew signal output
rlabel metal2 s 448610 0 448666 800 6 instrMgmt_dataOut[59]
port 158 nsew signal output
rlabel metal2 s 384026 0 384082 800 6 instrMgmt_dataOut[5]
port 159 nsew signal output
rlabel metal2 s 449806 0 449862 800 6 instrMgmt_dataOut[60]
port 160 nsew signal output
rlabel metal2 s 451002 0 451058 800 6 instrMgmt_dataOut[61]
port 161 nsew signal output
rlabel metal2 s 452198 0 452254 800 6 instrMgmt_dataOut[62]
port 162 nsew signal output
rlabel metal2 s 453394 0 453450 800 6 instrMgmt_dataOut[63]
port 163 nsew signal output
rlabel metal2 s 385222 0 385278 800 6 instrMgmt_dataOut[6]
port 164 nsew signal output
rlabel metal2 s 386418 0 386474 800 6 instrMgmt_dataOut[7]
port 165 nsew signal output
rlabel metal2 s 387614 0 387670 800 6 instrMgmt_dataOut[8]
port 166 nsew signal output
rlabel metal2 s 388810 0 388866 800 6 instrMgmt_dataOut[9]
port 167 nsew signal output
rlabel metal2 s 455786 0 455842 800 6 instrMgmt_we
port 168 nsew signal output
rlabel metal2 s 456982 0 457038 800 6 instrMgmt_wm[0]
port 169 nsew signal output
rlabel metal2 s 458178 0 458234 800 6 instrMgmt_wm[1]
port 170 nsew signal output
rlabel metal2 s 459374 0 459430 800 6 instrMgmt_wm[2]
port 171 nsew signal output
rlabel metal2 s 460570 0 460626 800 6 instrMgmt_wm[3]
port 172 nsew signal output
rlabel metal2 s 461766 0 461822 800 6 instrMgmt_wm[4]
port 173 nsew signal output
rlabel metal2 s 462962 0 463018 800 6 instrMgmt_wm[5]
port 174 nsew signal output
rlabel metal2 s 464158 0 464214 800 6 instrMgmt_wm[6]
port 175 nsew signal output
rlabel metal2 s 465354 0 465410 800 6 instrMgmt_wm[7]
port 176 nsew signal output
rlabel metal2 s 466550 0 466606 800 6 instr_addr[0]
port 177 nsew signal output
rlabel metal2 s 467746 0 467802 800 6 instr_addr[1]
port 178 nsew signal output
rlabel metal2 s 468942 0 468998 800 6 instr_addr[2]
port 179 nsew signal output
rlabel metal2 s 470138 0 470194 800 6 instr_addr[3]
port 180 nsew signal output
rlabel metal2 s 471334 0 471390 800 6 instr_addr[4]
port 181 nsew signal output
rlabel metal2 s 472530 0 472586 800 6 instr_addr[5]
port 182 nsew signal output
rlabel metal2 s 473726 0 473782 800 6 instr_addr[6]
port 183 nsew signal output
rlabel metal2 s 474922 0 474978 800 6 instr_addr[7]
port 184 nsew signal output
rlabel metal2 s 476118 0 476174 800 6 instr_addr[8]
port 185 nsew signal output
rlabel metal2 s 553858 0 553914 800 6 instr_ce
port 186 nsew signal output
rlabel metal2 s 477314 0 477370 800 6 instr_dataIn[0]
port 187 nsew signal input
rlabel metal2 s 489274 0 489330 800 6 instr_dataIn[10]
port 188 nsew signal input
rlabel metal2 s 490470 0 490526 800 6 instr_dataIn[11]
port 189 nsew signal input
rlabel metal2 s 491666 0 491722 800 6 instr_dataIn[12]
port 190 nsew signal input
rlabel metal2 s 492862 0 492918 800 6 instr_dataIn[13]
port 191 nsew signal input
rlabel metal2 s 494058 0 494114 800 6 instr_dataIn[14]
port 192 nsew signal input
rlabel metal2 s 495254 0 495310 800 6 instr_dataIn[15]
port 193 nsew signal input
rlabel metal2 s 496450 0 496506 800 6 instr_dataIn[16]
port 194 nsew signal input
rlabel metal2 s 497646 0 497702 800 6 instr_dataIn[17]
port 195 nsew signal input
rlabel metal2 s 498842 0 498898 800 6 instr_dataIn[18]
port 196 nsew signal input
rlabel metal2 s 500038 0 500094 800 6 instr_dataIn[19]
port 197 nsew signal input
rlabel metal2 s 478510 0 478566 800 6 instr_dataIn[1]
port 198 nsew signal input
rlabel metal2 s 501234 0 501290 800 6 instr_dataIn[20]
port 199 nsew signal input
rlabel metal2 s 502430 0 502486 800 6 instr_dataIn[21]
port 200 nsew signal input
rlabel metal2 s 503626 0 503682 800 6 instr_dataIn[22]
port 201 nsew signal input
rlabel metal2 s 504822 0 504878 800 6 instr_dataIn[23]
port 202 nsew signal input
rlabel metal2 s 506018 0 506074 800 6 instr_dataIn[24]
port 203 nsew signal input
rlabel metal2 s 507214 0 507270 800 6 instr_dataIn[25]
port 204 nsew signal input
rlabel metal2 s 508410 0 508466 800 6 instr_dataIn[26]
port 205 nsew signal input
rlabel metal2 s 509606 0 509662 800 6 instr_dataIn[27]
port 206 nsew signal input
rlabel metal2 s 510802 0 510858 800 6 instr_dataIn[28]
port 207 nsew signal input
rlabel metal2 s 511998 0 512054 800 6 instr_dataIn[29]
port 208 nsew signal input
rlabel metal2 s 479706 0 479762 800 6 instr_dataIn[2]
port 209 nsew signal input
rlabel metal2 s 513194 0 513250 800 6 instr_dataIn[30]
port 210 nsew signal input
rlabel metal2 s 514390 0 514446 800 6 instr_dataIn[31]
port 211 nsew signal input
rlabel metal2 s 515586 0 515642 800 6 instr_dataIn[32]
port 212 nsew signal input
rlabel metal2 s 516782 0 516838 800 6 instr_dataIn[33]
port 213 nsew signal input
rlabel metal2 s 517978 0 518034 800 6 instr_dataIn[34]
port 214 nsew signal input
rlabel metal2 s 519174 0 519230 800 6 instr_dataIn[35]
port 215 nsew signal input
rlabel metal2 s 520370 0 520426 800 6 instr_dataIn[36]
port 216 nsew signal input
rlabel metal2 s 521566 0 521622 800 6 instr_dataIn[37]
port 217 nsew signal input
rlabel metal2 s 522762 0 522818 800 6 instr_dataIn[38]
port 218 nsew signal input
rlabel metal2 s 523958 0 524014 800 6 instr_dataIn[39]
port 219 nsew signal input
rlabel metal2 s 480902 0 480958 800 6 instr_dataIn[3]
port 220 nsew signal input
rlabel metal2 s 525154 0 525210 800 6 instr_dataIn[40]
port 221 nsew signal input
rlabel metal2 s 526350 0 526406 800 6 instr_dataIn[41]
port 222 nsew signal input
rlabel metal2 s 527546 0 527602 800 6 instr_dataIn[42]
port 223 nsew signal input
rlabel metal2 s 528742 0 528798 800 6 instr_dataIn[43]
port 224 nsew signal input
rlabel metal2 s 529938 0 529994 800 6 instr_dataIn[44]
port 225 nsew signal input
rlabel metal2 s 531134 0 531190 800 6 instr_dataIn[45]
port 226 nsew signal input
rlabel metal2 s 532330 0 532386 800 6 instr_dataIn[46]
port 227 nsew signal input
rlabel metal2 s 533526 0 533582 800 6 instr_dataIn[47]
port 228 nsew signal input
rlabel metal2 s 534722 0 534778 800 6 instr_dataIn[48]
port 229 nsew signal input
rlabel metal2 s 535918 0 535974 800 6 instr_dataIn[49]
port 230 nsew signal input
rlabel metal2 s 482098 0 482154 800 6 instr_dataIn[4]
port 231 nsew signal input
rlabel metal2 s 537114 0 537170 800 6 instr_dataIn[50]
port 232 nsew signal input
rlabel metal2 s 538310 0 538366 800 6 instr_dataIn[51]
port 233 nsew signal input
rlabel metal2 s 539506 0 539562 800 6 instr_dataIn[52]
port 234 nsew signal input
rlabel metal2 s 540702 0 540758 800 6 instr_dataIn[53]
port 235 nsew signal input
rlabel metal2 s 541898 0 541954 800 6 instr_dataIn[54]
port 236 nsew signal input
rlabel metal2 s 543094 0 543150 800 6 instr_dataIn[55]
port 237 nsew signal input
rlabel metal2 s 544290 0 544346 800 6 instr_dataIn[56]
port 238 nsew signal input
rlabel metal2 s 545486 0 545542 800 6 instr_dataIn[57]
port 239 nsew signal input
rlabel metal2 s 546682 0 546738 800 6 instr_dataIn[58]
port 240 nsew signal input
rlabel metal2 s 547878 0 547934 800 6 instr_dataIn[59]
port 241 nsew signal input
rlabel metal2 s 483294 0 483350 800 6 instr_dataIn[5]
port 242 nsew signal input
rlabel metal2 s 549074 0 549130 800 6 instr_dataIn[60]
port 243 nsew signal input
rlabel metal2 s 550270 0 550326 800 6 instr_dataIn[61]
port 244 nsew signal input
rlabel metal2 s 551466 0 551522 800 6 instr_dataIn[62]
port 245 nsew signal input
rlabel metal2 s 552662 0 552718 800 6 instr_dataIn[63]
port 246 nsew signal input
rlabel metal2 s 484490 0 484546 800 6 instr_dataIn[6]
port 247 nsew signal input
rlabel metal2 s 485686 0 485742 800 6 instr_dataIn[7]
port 248 nsew signal input
rlabel metal2 s 486882 0 486938 800 6 instr_dataIn[8]
port 249 nsew signal input
rlabel metal2 s 488078 0 488134 800 6 instr_dataIn[9]
port 250 nsew signal input
rlabel metal3 s 559200 5856 560000 5976 6 io_in[0]
port 251 nsew signal input
rlabel metal3 s 559200 287376 560000 287496 6 io_in[10]
port 252 nsew signal input
rlabel metal3 s 559200 315528 560000 315648 6 io_in[11]
port 253 nsew signal input
rlabel metal3 s 559200 343680 560000 343800 6 io_in[12]
port 254 nsew signal input
rlabel metal3 s 559200 371832 560000 371952 6 io_in[13]
port 255 nsew signal input
rlabel metal3 s 559200 399984 560000 400104 6 io_in[14]
port 256 nsew signal input
rlabel metal2 s 430670 499200 430726 500000 6 io_in[15]
port 257 nsew signal input
rlabel metal2 s 445022 499200 445078 500000 6 io_in[16]
port 258 nsew signal input
rlabel metal2 s 459374 499200 459430 500000 6 io_in[17]
port 259 nsew signal input
rlabel metal2 s 473726 499200 473782 500000 6 io_in[18]
port 260 nsew signal input
rlabel metal2 s 488078 499200 488134 500000 6 io_in[19]
port 261 nsew signal input
rlabel metal3 s 559200 34008 560000 34128 6 io_in[1]
port 262 nsew signal input
rlabel metal2 s 502430 499200 502486 500000 6 io_in[20]
port 263 nsew signal input
rlabel metal2 s 516782 499200 516838 500000 6 io_in[21]
port 264 nsew signal input
rlabel metal2 s 531134 499200 531190 500000 6 io_in[22]
port 265 nsew signal input
rlabel metal2 s 545486 499200 545542 500000 6 io_in[23]
port 266 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[24]
port 267 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 io_in[25]
port 268 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 io_in[26]
port 269 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 io_in[27]
port 270 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 io_in[28]
port 271 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 io_in[29]
port 272 nsew signal input
rlabel metal3 s 559200 62160 560000 62280 6 io_in[2]
port 273 nsew signal input
rlabel metal3 s 0 171232 800 171352 6 io_in[30]
port 274 nsew signal input
rlabel metal3 s 0 198976 800 199096 6 io_in[31]
port 275 nsew signal input
rlabel metal3 s 0 226720 800 226840 6 io_in[32]
port 276 nsew signal input
rlabel metal3 s 0 254464 800 254584 6 io_in[33]
port 277 nsew signal input
rlabel metal3 s 0 282208 800 282328 6 io_in[34]
port 278 nsew signal input
rlabel metal3 s 0 309952 800 310072 6 io_in[35]
port 279 nsew signal input
rlabel metal3 s 0 337696 800 337816 6 io_in[36]
port 280 nsew signal input
rlabel metal3 s 0 365440 800 365560 6 io_in[37]
port 281 nsew signal input
rlabel metal3 s 559200 90312 560000 90432 6 io_in[3]
port 282 nsew signal input
rlabel metal3 s 559200 118464 560000 118584 6 io_in[4]
port 283 nsew signal input
rlabel metal3 s 559200 146616 560000 146736 6 io_in[5]
port 284 nsew signal input
rlabel metal3 s 559200 174768 560000 174888 6 io_in[6]
port 285 nsew signal input
rlabel metal3 s 559200 202920 560000 203040 6 io_in[7]
port 286 nsew signal input
rlabel metal3 s 559200 231072 560000 231192 6 io_in[8]
port 287 nsew signal input
rlabel metal3 s 559200 259224 560000 259344 6 io_in[9]
port 288 nsew signal input
rlabel metal3 s 559200 15240 560000 15360 6 io_oeb[0]
port 289 nsew signal output
rlabel metal3 s 559200 296760 560000 296880 6 io_oeb[10]
port 290 nsew signal output
rlabel metal3 s 559200 324912 560000 325032 6 io_oeb[11]
port 291 nsew signal output
rlabel metal3 s 559200 353064 560000 353184 6 io_oeb[12]
port 292 nsew signal output
rlabel metal3 s 559200 381216 560000 381336 6 io_oeb[13]
port 293 nsew signal output
rlabel metal3 s 559200 409368 560000 409488 6 io_oeb[14]
port 294 nsew signal output
rlabel metal2 s 435454 499200 435510 500000 6 io_oeb[15]
port 295 nsew signal output
rlabel metal2 s 449806 499200 449862 500000 6 io_oeb[16]
port 296 nsew signal output
rlabel metal2 s 464158 499200 464214 500000 6 io_oeb[17]
port 297 nsew signal output
rlabel metal2 s 478510 499200 478566 500000 6 io_oeb[18]
port 298 nsew signal output
rlabel metal2 s 492862 499200 492918 500000 6 io_oeb[19]
port 299 nsew signal output
rlabel metal3 s 559200 43392 560000 43512 6 io_oeb[1]
port 300 nsew signal output
rlabel metal2 s 507214 499200 507270 500000 6 io_oeb[20]
port 301 nsew signal output
rlabel metal2 s 521566 499200 521622 500000 6 io_oeb[21]
port 302 nsew signal output
rlabel metal2 s 535918 499200 535974 500000 6 io_oeb[22]
port 303 nsew signal output
rlabel metal2 s 550270 499200 550326 500000 6 io_oeb[23]
port 304 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_oeb[24]
port 305 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 io_oeb[25]
port 306 nsew signal output
rlabel metal3 s 0 69504 800 69624 6 io_oeb[26]
port 307 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 io_oeb[27]
port 308 nsew signal output
rlabel metal3 s 0 124992 800 125112 6 io_oeb[28]
port 309 nsew signal output
rlabel metal3 s 0 152736 800 152856 6 io_oeb[29]
port 310 nsew signal output
rlabel metal3 s 559200 71544 560000 71664 6 io_oeb[2]
port 311 nsew signal output
rlabel metal3 s 0 180480 800 180600 6 io_oeb[30]
port 312 nsew signal output
rlabel metal3 s 0 208224 800 208344 6 io_oeb[31]
port 313 nsew signal output
rlabel metal3 s 0 235968 800 236088 6 io_oeb[32]
port 314 nsew signal output
rlabel metal3 s 0 263712 800 263832 6 io_oeb[33]
port 315 nsew signal output
rlabel metal3 s 0 291456 800 291576 6 io_oeb[34]
port 316 nsew signal output
rlabel metal3 s 0 319200 800 319320 6 io_oeb[35]
port 317 nsew signal output
rlabel metal3 s 0 346944 800 347064 6 io_oeb[36]
port 318 nsew signal output
rlabel metal3 s 0 374688 800 374808 6 io_oeb[37]
port 319 nsew signal output
rlabel metal3 s 559200 99696 560000 99816 6 io_oeb[3]
port 320 nsew signal output
rlabel metal3 s 559200 127848 560000 127968 6 io_oeb[4]
port 321 nsew signal output
rlabel metal3 s 559200 156000 560000 156120 6 io_oeb[5]
port 322 nsew signal output
rlabel metal3 s 559200 184152 560000 184272 6 io_oeb[6]
port 323 nsew signal output
rlabel metal3 s 559200 212304 560000 212424 6 io_oeb[7]
port 324 nsew signal output
rlabel metal3 s 559200 240456 560000 240576 6 io_oeb[8]
port 325 nsew signal output
rlabel metal3 s 559200 268608 560000 268728 6 io_oeb[9]
port 326 nsew signal output
rlabel metal3 s 559200 24624 560000 24744 6 io_out[0]
port 327 nsew signal output
rlabel metal3 s 559200 306144 560000 306264 6 io_out[10]
port 328 nsew signal output
rlabel metal3 s 559200 334296 560000 334416 6 io_out[11]
port 329 nsew signal output
rlabel metal3 s 559200 362448 560000 362568 6 io_out[12]
port 330 nsew signal output
rlabel metal3 s 559200 390600 560000 390720 6 io_out[13]
port 331 nsew signal output
rlabel metal3 s 559200 418752 560000 418872 6 io_out[14]
port 332 nsew signal output
rlabel metal2 s 440238 499200 440294 500000 6 io_out[15]
port 333 nsew signal output
rlabel metal2 s 454590 499200 454646 500000 6 io_out[16]
port 334 nsew signal output
rlabel metal2 s 468942 499200 468998 500000 6 io_out[17]
port 335 nsew signal output
rlabel metal2 s 483294 499200 483350 500000 6 io_out[18]
port 336 nsew signal output
rlabel metal2 s 497646 499200 497702 500000 6 io_out[19]
port 337 nsew signal output
rlabel metal3 s 559200 52776 560000 52896 6 io_out[1]
port 338 nsew signal output
rlabel metal2 s 511998 499200 512054 500000 6 io_out[20]
port 339 nsew signal output
rlabel metal2 s 526350 499200 526406 500000 6 io_out[21]
port 340 nsew signal output
rlabel metal2 s 540702 499200 540758 500000 6 io_out[22]
port 341 nsew signal output
rlabel metal2 s 555054 499200 555110 500000 6 io_out[23]
port 342 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 io_out[24]
port 343 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_out[25]
port 344 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 io_out[26]
port 345 nsew signal output
rlabel metal3 s 0 106496 800 106616 6 io_out[27]
port 346 nsew signal output
rlabel metal3 s 0 134240 800 134360 6 io_out[28]
port 347 nsew signal output
rlabel metal3 s 0 161984 800 162104 6 io_out[29]
port 348 nsew signal output
rlabel metal3 s 559200 80928 560000 81048 6 io_out[2]
port 349 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 io_out[30]
port 350 nsew signal output
rlabel metal3 s 0 217472 800 217592 6 io_out[31]
port 351 nsew signal output
rlabel metal3 s 0 245216 800 245336 6 io_out[32]
port 352 nsew signal output
rlabel metal3 s 0 272960 800 273080 6 io_out[33]
port 353 nsew signal output
rlabel metal3 s 0 300704 800 300824 6 io_out[34]
port 354 nsew signal output
rlabel metal3 s 0 328448 800 328568 6 io_out[35]
port 355 nsew signal output
rlabel metal3 s 0 356192 800 356312 6 io_out[36]
port 356 nsew signal output
rlabel metal3 s 0 383936 800 384056 6 io_out[37]
port 357 nsew signal output
rlabel metal3 s 559200 109080 560000 109200 6 io_out[3]
port 358 nsew signal output
rlabel metal3 s 559200 137232 560000 137352 6 io_out[4]
port 359 nsew signal output
rlabel metal3 s 559200 165384 560000 165504 6 io_out[5]
port 360 nsew signal output
rlabel metal3 s 559200 193536 560000 193656 6 io_out[6]
port 361 nsew signal output
rlabel metal3 s 559200 221688 560000 221808 6 io_out[7]
port 362 nsew signal output
rlabel metal3 s 559200 249840 560000 249960 6 io_out[8]
port 363 nsew signal output
rlabel metal3 s 559200 277992 560000 278112 6 io_out[9]
port 364 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 irq[0]
port 365 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 irq[1]
port 366 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 irq[2]
port 367 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[0]
port 368 nsew signal output
rlabel metal2 s 257250 0 257306 800 6 la_data_out[100]
port 369 nsew signal output
rlabel metal2 s 258446 0 258502 800 6 la_data_out[101]
port 370 nsew signal output
rlabel metal2 s 259642 0 259698 800 6 la_data_out[102]
port 371 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 la_data_out[103]
port 372 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 la_data_out[104]
port 373 nsew signal output
rlabel metal2 s 263230 0 263286 800 6 la_data_out[105]
port 374 nsew signal output
rlabel metal2 s 264426 0 264482 800 6 la_data_out[106]
port 375 nsew signal output
rlabel metal2 s 265622 0 265678 800 6 la_data_out[107]
port 376 nsew signal output
rlabel metal2 s 266818 0 266874 800 6 la_data_out[108]
port 377 nsew signal output
rlabel metal2 s 268014 0 268070 800 6 la_data_out[109]
port 378 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[10]
port 379 nsew signal output
rlabel metal2 s 269210 0 269266 800 6 la_data_out[110]
port 380 nsew signal output
rlabel metal2 s 270406 0 270462 800 6 la_data_out[111]
port 381 nsew signal output
rlabel metal2 s 271602 0 271658 800 6 la_data_out[112]
port 382 nsew signal output
rlabel metal2 s 272798 0 272854 800 6 la_data_out[113]
port 383 nsew signal output
rlabel metal2 s 273994 0 274050 800 6 la_data_out[114]
port 384 nsew signal output
rlabel metal2 s 275190 0 275246 800 6 la_data_out[115]
port 385 nsew signal output
rlabel metal2 s 276386 0 276442 800 6 la_data_out[116]
port 386 nsew signal output
rlabel metal2 s 277582 0 277638 800 6 la_data_out[117]
port 387 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[118]
port 388 nsew signal output
rlabel metal2 s 279974 0 280030 800 6 la_data_out[119]
port 389 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 la_data_out[11]
port 390 nsew signal output
rlabel metal2 s 281170 0 281226 800 6 la_data_out[120]
port 391 nsew signal output
rlabel metal2 s 282366 0 282422 800 6 la_data_out[121]
port 392 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 la_data_out[122]
port 393 nsew signal output
rlabel metal2 s 284758 0 284814 800 6 la_data_out[123]
port 394 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[124]
port 395 nsew signal output
rlabel metal2 s 287150 0 287206 800 6 la_data_out[125]
port 396 nsew signal output
rlabel metal2 s 288346 0 288402 800 6 la_data_out[126]
port 397 nsew signal output
rlabel metal2 s 289542 0 289598 800 6 la_data_out[127]
port 398 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[12]
port 399 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[13]
port 400 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[14]
port 401 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[15]
port 402 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 la_data_out[16]
port 403 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 la_data_out[17]
port 404 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[18]
port 405 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[19]
port 406 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[1]
port 407 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 la_data_out[20]
port 408 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 la_data_out[21]
port 409 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[22]
port 410 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[23]
port 411 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[24]
port 412 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[25]
port 413 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[26]
port 414 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[27]
port 415 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[28]
port 416 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[29]
port 417 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[2]
port 418 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[30]
port 419 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[31]
port 420 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[32]
port 421 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 la_data_out[33]
port 422 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[34]
port 423 nsew signal output
rlabel metal2 s 179510 0 179566 800 6 la_data_out[35]
port 424 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[36]
port 425 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 la_data_out[37]
port 426 nsew signal output
rlabel metal2 s 183098 0 183154 800 6 la_data_out[38]
port 427 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[39]
port 428 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[3]
port 429 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[40]
port 430 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[41]
port 431 nsew signal output
rlabel metal2 s 187882 0 187938 800 6 la_data_out[42]
port 432 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[43]
port 433 nsew signal output
rlabel metal2 s 190274 0 190330 800 6 la_data_out[44]
port 434 nsew signal output
rlabel metal2 s 191470 0 191526 800 6 la_data_out[45]
port 435 nsew signal output
rlabel metal2 s 192666 0 192722 800 6 la_data_out[46]
port 436 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 la_data_out[47]
port 437 nsew signal output
rlabel metal2 s 195058 0 195114 800 6 la_data_out[48]
port 438 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[49]
port 439 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[4]
port 440 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[50]
port 441 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[51]
port 442 nsew signal output
rlabel metal2 s 199842 0 199898 800 6 la_data_out[52]
port 443 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[53]
port 444 nsew signal output
rlabel metal2 s 202234 0 202290 800 6 la_data_out[54]
port 445 nsew signal output
rlabel metal2 s 203430 0 203486 800 6 la_data_out[55]
port 446 nsew signal output
rlabel metal2 s 204626 0 204682 800 6 la_data_out[56]
port 447 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[57]
port 448 nsew signal output
rlabel metal2 s 207018 0 207074 800 6 la_data_out[58]
port 449 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[59]
port 450 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[5]
port 451 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[60]
port 452 nsew signal output
rlabel metal2 s 210606 0 210662 800 6 la_data_out[61]
port 453 nsew signal output
rlabel metal2 s 211802 0 211858 800 6 la_data_out[62]
port 454 nsew signal output
rlabel metal2 s 212998 0 213054 800 6 la_data_out[63]
port 455 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[64]
port 456 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 la_data_out[65]
port 457 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[66]
port 458 nsew signal output
rlabel metal2 s 217782 0 217838 800 6 la_data_out[67]
port 459 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[68]
port 460 nsew signal output
rlabel metal2 s 220174 0 220230 800 6 la_data_out[69]
port 461 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[6]
port 462 nsew signal output
rlabel metal2 s 221370 0 221426 800 6 la_data_out[70]
port 463 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[71]
port 464 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[72]
port 465 nsew signal output
rlabel metal2 s 224958 0 225014 800 6 la_data_out[73]
port 466 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[74]
port 467 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[75]
port 468 nsew signal output
rlabel metal2 s 228546 0 228602 800 6 la_data_out[76]
port 469 nsew signal output
rlabel metal2 s 229742 0 229798 800 6 la_data_out[77]
port 470 nsew signal output
rlabel metal2 s 230938 0 230994 800 6 la_data_out[78]
port 471 nsew signal output
rlabel metal2 s 232134 0 232190 800 6 la_data_out[79]
port 472 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[7]
port 473 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[80]
port 474 nsew signal output
rlabel metal2 s 234526 0 234582 800 6 la_data_out[81]
port 475 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 la_data_out[82]
port 476 nsew signal output
rlabel metal2 s 236918 0 236974 800 6 la_data_out[83]
port 477 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[84]
port 478 nsew signal output
rlabel metal2 s 239310 0 239366 800 6 la_data_out[85]
port 479 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[86]
port 480 nsew signal output
rlabel metal2 s 241702 0 241758 800 6 la_data_out[87]
port 481 nsew signal output
rlabel metal2 s 242898 0 242954 800 6 la_data_out[88]
port 482 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[89]
port 483 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[8]
port 484 nsew signal output
rlabel metal2 s 245290 0 245346 800 6 la_data_out[90]
port 485 nsew signal output
rlabel metal2 s 246486 0 246542 800 6 la_data_out[91]
port 486 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[92]
port 487 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[93]
port 488 nsew signal output
rlabel metal2 s 250074 0 250130 800 6 la_data_out[94]
port 489 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 la_data_out[95]
port 490 nsew signal output
rlabel metal2 s 252466 0 252522 800 6 la_data_out[96]
port 491 nsew signal output
rlabel metal2 s 253662 0 253718 800 6 la_data_out[97]
port 492 nsew signal output
rlabel metal2 s 254858 0 254914 800 6 la_data_out[98]
port 493 nsew signal output
rlabel metal2 s 256054 0 256110 800 6 la_data_out[99]
port 494 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[9]
port 495 nsew signal output
rlabel metal2 s 4894 499200 4950 500000 6 mem_addr[0]
port 496 nsew signal output
rlabel metal2 s 9678 499200 9734 500000 6 mem_addr[1]
port 497 nsew signal output
rlabel metal2 s 14462 499200 14518 500000 6 mem_addr[2]
port 498 nsew signal output
rlabel metal2 s 19246 499200 19302 500000 6 mem_addr[3]
port 499 nsew signal output
rlabel metal2 s 24030 499200 24086 500000 6 mem_addr[4]
port 500 nsew signal output
rlabel metal2 s 28814 499200 28870 500000 6 mem_addr[5]
port 501 nsew signal output
rlabel metal2 s 33598 499200 33654 500000 6 mem_addr[6]
port 502 nsew signal output
rlabel metal2 s 38382 499200 38438 500000 6 mem_addr[7]
port 503 nsew signal output
rlabel metal2 s 43166 499200 43222 500000 6 mem_addr[8]
port 504 nsew signal output
rlabel metal2 s 378046 499200 378102 500000 6 mem_ce
port 505 nsew signal output
rlabel metal2 s 47950 499200 48006 500000 6 mem_dataIn[0]
port 506 nsew signal input
rlabel metal2 s 95790 499200 95846 500000 6 mem_dataIn[10]
port 507 nsew signal input
rlabel metal2 s 100574 499200 100630 500000 6 mem_dataIn[11]
port 508 nsew signal input
rlabel metal2 s 105358 499200 105414 500000 6 mem_dataIn[12]
port 509 nsew signal input
rlabel metal2 s 110142 499200 110198 500000 6 mem_dataIn[13]
port 510 nsew signal input
rlabel metal2 s 114926 499200 114982 500000 6 mem_dataIn[14]
port 511 nsew signal input
rlabel metal2 s 119710 499200 119766 500000 6 mem_dataIn[15]
port 512 nsew signal input
rlabel metal2 s 124494 499200 124550 500000 6 mem_dataIn[16]
port 513 nsew signal input
rlabel metal2 s 129278 499200 129334 500000 6 mem_dataIn[17]
port 514 nsew signal input
rlabel metal2 s 134062 499200 134118 500000 6 mem_dataIn[18]
port 515 nsew signal input
rlabel metal2 s 138846 499200 138902 500000 6 mem_dataIn[19]
port 516 nsew signal input
rlabel metal2 s 52734 499200 52790 500000 6 mem_dataIn[1]
port 517 nsew signal input
rlabel metal2 s 143630 499200 143686 500000 6 mem_dataIn[20]
port 518 nsew signal input
rlabel metal2 s 148414 499200 148470 500000 6 mem_dataIn[21]
port 519 nsew signal input
rlabel metal2 s 153198 499200 153254 500000 6 mem_dataIn[22]
port 520 nsew signal input
rlabel metal2 s 157982 499200 158038 500000 6 mem_dataIn[23]
port 521 nsew signal input
rlabel metal2 s 162766 499200 162822 500000 6 mem_dataIn[24]
port 522 nsew signal input
rlabel metal2 s 167550 499200 167606 500000 6 mem_dataIn[25]
port 523 nsew signal input
rlabel metal2 s 172334 499200 172390 500000 6 mem_dataIn[26]
port 524 nsew signal input
rlabel metal2 s 177118 499200 177174 500000 6 mem_dataIn[27]
port 525 nsew signal input
rlabel metal2 s 181902 499200 181958 500000 6 mem_dataIn[28]
port 526 nsew signal input
rlabel metal2 s 186686 499200 186742 500000 6 mem_dataIn[29]
port 527 nsew signal input
rlabel metal2 s 57518 499200 57574 500000 6 mem_dataIn[2]
port 528 nsew signal input
rlabel metal2 s 191470 499200 191526 500000 6 mem_dataIn[30]
port 529 nsew signal input
rlabel metal2 s 196254 499200 196310 500000 6 mem_dataIn[31]
port 530 nsew signal input
rlabel metal2 s 62302 499200 62358 500000 6 mem_dataIn[3]
port 531 nsew signal input
rlabel metal2 s 67086 499200 67142 500000 6 mem_dataIn[4]
port 532 nsew signal input
rlabel metal2 s 71870 499200 71926 500000 6 mem_dataIn[5]
port 533 nsew signal input
rlabel metal2 s 76654 499200 76710 500000 6 mem_dataIn[6]
port 534 nsew signal input
rlabel metal2 s 81438 499200 81494 500000 6 mem_dataIn[7]
port 535 nsew signal input
rlabel metal2 s 86222 499200 86278 500000 6 mem_dataIn[8]
port 536 nsew signal input
rlabel metal2 s 91006 499200 91062 500000 6 mem_dataIn[9]
port 537 nsew signal input
rlabel metal2 s 201038 499200 201094 500000 6 mem_dataOut[0]
port 538 nsew signal output
rlabel metal2 s 248878 499200 248934 500000 6 mem_dataOut[10]
port 539 nsew signal output
rlabel metal2 s 253662 499200 253718 500000 6 mem_dataOut[11]
port 540 nsew signal output
rlabel metal2 s 258446 499200 258502 500000 6 mem_dataOut[12]
port 541 nsew signal output
rlabel metal2 s 263230 499200 263286 500000 6 mem_dataOut[13]
port 542 nsew signal output
rlabel metal2 s 268014 499200 268070 500000 6 mem_dataOut[14]
port 543 nsew signal output
rlabel metal2 s 272798 499200 272854 500000 6 mem_dataOut[15]
port 544 nsew signal output
rlabel metal2 s 277582 499200 277638 500000 6 mem_dataOut[16]
port 545 nsew signal output
rlabel metal2 s 282366 499200 282422 500000 6 mem_dataOut[17]
port 546 nsew signal output
rlabel metal2 s 287150 499200 287206 500000 6 mem_dataOut[18]
port 547 nsew signal output
rlabel metal2 s 291934 499200 291990 500000 6 mem_dataOut[19]
port 548 nsew signal output
rlabel metal2 s 205822 499200 205878 500000 6 mem_dataOut[1]
port 549 nsew signal output
rlabel metal2 s 296718 499200 296774 500000 6 mem_dataOut[20]
port 550 nsew signal output
rlabel metal2 s 301502 499200 301558 500000 6 mem_dataOut[21]
port 551 nsew signal output
rlabel metal2 s 306286 499200 306342 500000 6 mem_dataOut[22]
port 552 nsew signal output
rlabel metal2 s 311070 499200 311126 500000 6 mem_dataOut[23]
port 553 nsew signal output
rlabel metal2 s 315854 499200 315910 500000 6 mem_dataOut[24]
port 554 nsew signal output
rlabel metal2 s 320638 499200 320694 500000 6 mem_dataOut[25]
port 555 nsew signal output
rlabel metal2 s 325422 499200 325478 500000 6 mem_dataOut[26]
port 556 nsew signal output
rlabel metal2 s 330206 499200 330262 500000 6 mem_dataOut[27]
port 557 nsew signal output
rlabel metal2 s 334990 499200 335046 500000 6 mem_dataOut[28]
port 558 nsew signal output
rlabel metal2 s 339774 499200 339830 500000 6 mem_dataOut[29]
port 559 nsew signal output
rlabel metal2 s 210606 499200 210662 500000 6 mem_dataOut[2]
port 560 nsew signal output
rlabel metal2 s 344558 499200 344614 500000 6 mem_dataOut[30]
port 561 nsew signal output
rlabel metal2 s 349342 499200 349398 500000 6 mem_dataOut[31]
port 562 nsew signal output
rlabel metal2 s 215390 499200 215446 500000 6 mem_dataOut[3]
port 563 nsew signal output
rlabel metal2 s 220174 499200 220230 500000 6 mem_dataOut[4]
port 564 nsew signal output
rlabel metal2 s 224958 499200 225014 500000 6 mem_dataOut[5]
port 565 nsew signal output
rlabel metal2 s 229742 499200 229798 500000 6 mem_dataOut[6]
port 566 nsew signal output
rlabel metal2 s 234526 499200 234582 500000 6 mem_dataOut[7]
port 567 nsew signal output
rlabel metal2 s 239310 499200 239366 500000 6 mem_dataOut[8]
port 568 nsew signal output
rlabel metal2 s 244094 499200 244150 500000 6 mem_dataOut[9]
port 569 nsew signal output
rlabel metal2 s 373262 499200 373318 500000 6 mem_we
port 570 nsew signal output
rlabel metal2 s 354126 499200 354182 500000 6 mem_wm[0]
port 571 nsew signal output
rlabel metal2 s 358910 499200 358966 500000 6 mem_wm[1]
port 572 nsew signal output
rlabel metal2 s 363694 499200 363750 500000 6 mem_wm[2]
port 573 nsew signal output
rlabel metal2 s 368478 499200 368534 500000 6 mem_wm[3]
port 574 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 user_clock2
port 575 nsew signal input
rlabel metal4 s 4208 2128 4528 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 497808 6 vccd1
port 576 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 497808 6 vssd1
port 577 nsew ground bidirectional
rlabel metal2 s 135258 0 135314 800 6 wb_clk_i
port 578 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 wb_rst_i
port 579 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_ack_o
port 580 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[0]
port 581 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_adr_i[10]
port 582 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_adr_i[11]
port 583 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_adr_i[12]
port 584 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 wbs_adr_i[13]
port 585 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 wbs_adr_i[14]
port 586 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_adr_i[15]
port 587 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_adr_i[16]
port 588 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wbs_adr_i[17]
port 589 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_adr_i[18]
port 590 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 wbs_adr_i[19]
port 591 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[1]
port 592 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 wbs_adr_i[20]
port 593 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 wbs_adr_i[21]
port 594 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 wbs_adr_i[22]
port 595 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 wbs_adr_i[23]
port 596 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 wbs_adr_i[24]
port 597 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 wbs_adr_i[25]
port 598 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wbs_adr_i[26]
port 599 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 wbs_adr_i[27]
port 600 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 wbs_adr_i[28]
port 601 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 wbs_adr_i[29]
port 602 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_adr_i[2]
port 603 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 wbs_adr_i[30]
port 604 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 wbs_adr_i[31]
port 605 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[3]
port 606 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[4]
port 607 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_adr_i[5]
port 608 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[6]
port 609 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_adr_i[7]
port 610 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_adr_i[8]
port 611 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[9]
port 612 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_cyc_i
port 613 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 wbs_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 wbs_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 wbs_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 wbs_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 wbs_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 wbs_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 wbs_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 wbs_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 wbs_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 wbs_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[0]
port 646 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[10]
port 647 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[11]
port 648 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_o[12]
port 649 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_o[13]
port 650 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 wbs_dat_o[14]
port 651 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_o[15]
port 652 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 wbs_dat_o[16]
port 653 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 wbs_dat_o[17]
port 654 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[18]
port 655 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 wbs_dat_o[19]
port 656 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[1]
port 657 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 wbs_dat_o[20]
port 658 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_o[21]
port 659 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_o[22]
port 660 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 wbs_dat_o[23]
port 661 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 wbs_dat_o[24]
port 662 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 wbs_dat_o[25]
port 663 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 wbs_dat_o[26]
port 664 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 wbs_dat_o[27]
port 665 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 wbs_dat_o[28]
port 666 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 wbs_dat_o[29]
port 667 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[2]
port 668 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 wbs_dat_o[30]
port 669 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 wbs_dat_o[31]
port 670 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[3]
port 671 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_o[4]
port 672 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_o[5]
port 673 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[6]
port 674 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_o[7]
port 675 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[8]
port 676 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_o[9]
port 677 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_sel_i[0]
port 678 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_sel_i[1]
port 679 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_sel_i[2]
port 680 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_sel_i[3]
port 681 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_stb_i
port 682 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_we_i
port 683 nsew signal input
rlabel metal2 s 382830 499200 382886 500000 6 zero
port 684 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 560000 500000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 551601486
string GDS_FILE /home/m/Builds/Caraval/openlane/soomrv/runs/22_09_11_14_56/results/signoff/soomrv.magic.gds
string GDS_START 2069086
<< end >>

