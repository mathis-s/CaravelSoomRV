VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO soomrv
  CLASS BLOCK ;
  FOREIGN soomrv ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 2500.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2140.680 2800.000 2141.280 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 2496.000 1986.190 2500.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.830 2496.000 2010.110 2500.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.750 2496.000 2034.030 2500.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 2496.000 2057.950 2500.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.590 2496.000 2081.870 2500.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.510 2496.000 2105.790 2500.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.430 2496.000 2129.710 2500.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1965.920 4.000 1966.520 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.160 4.000 2012.760 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2058.400 4.000 2059.000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2187.600 2800.000 2188.200 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2104.640 4.000 2105.240 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2150.880 4.000 2151.480 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2197.120 4.000 2197.720 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2243.360 4.000 2243.960 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2289.600 4.000 2290.200 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2335.840 4.000 2336.440 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2382.080 4.000 2382.680 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2428.320 4.000 2428.920 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2474.560 4.000 2475.160 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2234.520 2800.000 2235.120 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2281.440 2800.000 2282.040 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2328.360 2800.000 2328.960 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2375.280 2800.000 2375.880 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2422.200 2800.000 2422.800 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2469.120 2800.000 2469.720 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 2496.000 1938.350 2500.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.990 2496.000 1962.270 2500.000 ;
    END
  END analog_io[9]
  PIN instrMgmt_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END instrMgmt_addr[0]
  PIN instrMgmt_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 0.000 1459.950 4.000 ;
    END
  END instrMgmt_addr[1]
  PIN instrMgmt_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.650 0.000 1465.930 4.000 ;
    END
  END instrMgmt_addr[2]
  PIN instrMgmt_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END instrMgmt_addr[3]
  PIN instrMgmt_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 0.000 1477.890 4.000 ;
    END
  END instrMgmt_addr[4]
  PIN instrMgmt_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 0.000 1483.870 4.000 ;
    END
  END instrMgmt_addr[5]
  PIN instrMgmt_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.570 0.000 1489.850 4.000 ;
    END
  END instrMgmt_addr[6]
  PIN instrMgmt_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END instrMgmt_addr[7]
  PIN instrMgmt_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END instrMgmt_addr[8]
  PIN instrMgmt_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.950 0.000 2273.230 4.000 ;
    END
  END instrMgmt_ce
  PIN instrMgmt_dataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 0.000 1507.790 4.000 ;
    END
  END instrMgmt_dataIn[0]
  PIN instrMgmt_dataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 0.000 1567.590 4.000 ;
    END
  END instrMgmt_dataIn[10]
  PIN instrMgmt_dataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 0.000 1573.570 4.000 ;
    END
  END instrMgmt_dataIn[11]
  PIN instrMgmt_dataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 0.000 1579.550 4.000 ;
    END
  END instrMgmt_dataIn[12]
  PIN instrMgmt_dataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.250 0.000 1585.530 4.000 ;
    END
  END instrMgmt_dataIn[13]
  PIN instrMgmt_dataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 0.000 1591.510 4.000 ;
    END
  END instrMgmt_dataIn[14]
  PIN instrMgmt_dataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END instrMgmt_dataIn[15]
  PIN instrMgmt_dataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.190 0.000 1603.470 4.000 ;
    END
  END instrMgmt_dataIn[16]
  PIN instrMgmt_dataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 0.000 1609.450 4.000 ;
    END
  END instrMgmt_dataIn[17]
  PIN instrMgmt_dataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END instrMgmt_dataIn[18]
  PIN instrMgmt_dataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 0.000 1621.410 4.000 ;
    END
  END instrMgmt_dataIn[19]
  PIN instrMgmt_dataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END instrMgmt_dataIn[1]
  PIN instrMgmt_dataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 0.000 1627.390 4.000 ;
    END
  END instrMgmt_dataIn[20]
  PIN instrMgmt_dataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 0.000 1633.370 4.000 ;
    END
  END instrMgmt_dataIn[21]
  PIN instrMgmt_dataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 0.000 1639.350 4.000 ;
    END
  END instrMgmt_dataIn[22]
  PIN instrMgmt_dataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 0.000 1645.330 4.000 ;
    END
  END instrMgmt_dataIn[23]
  PIN instrMgmt_dataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 0.000 1651.310 4.000 ;
    END
  END instrMgmt_dataIn[24]
  PIN instrMgmt_dataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.010 0.000 1657.290 4.000 ;
    END
  END instrMgmt_dataIn[25]
  PIN instrMgmt_dataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 0.000 1663.270 4.000 ;
    END
  END instrMgmt_dataIn[26]
  PIN instrMgmt_dataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 0.000 1669.250 4.000 ;
    END
  END instrMgmt_dataIn[27]
  PIN instrMgmt_dataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 0.000 1675.230 4.000 ;
    END
  END instrMgmt_dataIn[28]
  PIN instrMgmt_dataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END instrMgmt_dataIn[29]
  PIN instrMgmt_dataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 0.000 1519.750 4.000 ;
    END
  END instrMgmt_dataIn[2]
  PIN instrMgmt_dataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 0.000 1687.190 4.000 ;
    END
  END instrMgmt_dataIn[30]
  PIN instrMgmt_dataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.890 0.000 1693.170 4.000 ;
    END
  END instrMgmt_dataIn[31]
  PIN instrMgmt_dataIn[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 0.000 1699.150 4.000 ;
    END
  END instrMgmt_dataIn[32]
  PIN instrMgmt_dataIn[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END instrMgmt_dataIn[33]
  PIN instrMgmt_dataIn[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.830 0.000 1711.110 4.000 ;
    END
  END instrMgmt_dataIn[34]
  PIN instrMgmt_dataIn[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 4.000 ;
    END
  END instrMgmt_dataIn[35]
  PIN instrMgmt_dataIn[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 0.000 1723.070 4.000 ;
    END
  END instrMgmt_dataIn[36]
  PIN instrMgmt_dataIn[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 0.000 1729.050 4.000 ;
    END
  END instrMgmt_dataIn[37]
  PIN instrMgmt_dataIn[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 0.000 1735.030 4.000 ;
    END
  END instrMgmt_dataIn[38]
  PIN instrMgmt_dataIn[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.730 0.000 1741.010 4.000 ;
    END
  END instrMgmt_dataIn[39]
  PIN instrMgmt_dataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.450 0.000 1525.730 4.000 ;
    END
  END instrMgmt_dataIn[3]
  PIN instrMgmt_dataIn[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.710 0.000 1746.990 4.000 ;
    END
  END instrMgmt_dataIn[40]
  PIN instrMgmt_dataIn[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 0.000 1752.970 4.000 ;
    END
  END instrMgmt_dataIn[41]
  PIN instrMgmt_dataIn[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.670 0.000 1758.950 4.000 ;
    END
  END instrMgmt_dataIn[42]
  PIN instrMgmt_dataIn[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 0.000 1764.930 4.000 ;
    END
  END instrMgmt_dataIn[43]
  PIN instrMgmt_dataIn[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 0.000 1770.910 4.000 ;
    END
  END instrMgmt_dataIn[44]
  PIN instrMgmt_dataIn[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.610 0.000 1776.890 4.000 ;
    END
  END instrMgmt_dataIn[45]
  PIN instrMgmt_dataIn[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.590 0.000 1782.870 4.000 ;
    END
  END instrMgmt_dataIn[46]
  PIN instrMgmt_dataIn[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.570 0.000 1788.850 4.000 ;
    END
  END instrMgmt_dataIn[47]
  PIN instrMgmt_dataIn[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.550 0.000 1794.830 4.000 ;
    END
  END instrMgmt_dataIn[48]
  PIN instrMgmt_dataIn[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 0.000 1800.810 4.000 ;
    END
  END instrMgmt_dataIn[49]
  PIN instrMgmt_dataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.430 0.000 1531.710 4.000 ;
    END
  END instrMgmt_dataIn[4]
  PIN instrMgmt_dataIn[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END instrMgmt_dataIn[50]
  PIN instrMgmt_dataIn[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.490 0.000 1812.770 4.000 ;
    END
  END instrMgmt_dataIn[51]
  PIN instrMgmt_dataIn[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.470 0.000 1818.750 4.000 ;
    END
  END instrMgmt_dataIn[52]
  PIN instrMgmt_dataIn[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.450 0.000 1824.730 4.000 ;
    END
  END instrMgmt_dataIn[53]
  PIN instrMgmt_dataIn[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.430 0.000 1830.710 4.000 ;
    END
  END instrMgmt_dataIn[54]
  PIN instrMgmt_dataIn[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.410 0.000 1836.690 4.000 ;
    END
  END instrMgmt_dataIn[55]
  PIN instrMgmt_dataIn[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.390 0.000 1842.670 4.000 ;
    END
  END instrMgmt_dataIn[56]
  PIN instrMgmt_dataIn[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 0.000 1848.650 4.000 ;
    END
  END instrMgmt_dataIn[57]
  PIN instrMgmt_dataIn[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.350 0.000 1854.630 4.000 ;
    END
  END instrMgmt_dataIn[58]
  PIN instrMgmt_dataIn[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.330 0.000 1860.610 4.000 ;
    END
  END instrMgmt_dataIn[59]
  PIN instrMgmt_dataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 0.000 1537.690 4.000 ;
    END
  END instrMgmt_dataIn[5]
  PIN instrMgmt_dataIn[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.310 0.000 1866.590 4.000 ;
    END
  END instrMgmt_dataIn[60]
  PIN instrMgmt_dataIn[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.290 0.000 1872.570 4.000 ;
    END
  END instrMgmt_dataIn[61]
  PIN instrMgmt_dataIn[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.270 0.000 1878.550 4.000 ;
    END
  END instrMgmt_dataIn[62]
  PIN instrMgmt_dataIn[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.250 0.000 1884.530 4.000 ;
    END
  END instrMgmt_dataIn[63]
  PIN instrMgmt_dataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.390 0.000 1543.670 4.000 ;
    END
  END instrMgmt_dataIn[6]
  PIN instrMgmt_dataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.370 0.000 1549.650 4.000 ;
    END
  END instrMgmt_dataIn[7]
  PIN instrMgmt_dataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END instrMgmt_dataIn[8]
  PIN instrMgmt_dataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 0.000 1561.610 4.000 ;
    END
  END instrMgmt_dataIn[9]
  PIN instrMgmt_dataOut[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 0.000 1890.510 4.000 ;
    END
  END instrMgmt_dataOut[0]
  PIN instrMgmt_dataOut[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 0.000 1950.310 4.000 ;
    END
  END instrMgmt_dataOut[10]
  PIN instrMgmt_dataOut[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END instrMgmt_dataOut[11]
  PIN instrMgmt_dataOut[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.990 0.000 1962.270 4.000 ;
    END
  END instrMgmt_dataOut[12]
  PIN instrMgmt_dataOut[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.970 0.000 1968.250 4.000 ;
    END
  END instrMgmt_dataOut[13]
  PIN instrMgmt_dataOut[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 0.000 1974.230 4.000 ;
    END
  END instrMgmt_dataOut[14]
  PIN instrMgmt_dataOut[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.930 0.000 1980.210 4.000 ;
    END
  END instrMgmt_dataOut[15]
  PIN instrMgmt_dataOut[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 0.000 1986.190 4.000 ;
    END
  END instrMgmt_dataOut[16]
  PIN instrMgmt_dataOut[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.890 0.000 1992.170 4.000 ;
    END
  END instrMgmt_dataOut[17]
  PIN instrMgmt_dataOut[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.870 0.000 1998.150 4.000 ;
    END
  END instrMgmt_dataOut[18]
  PIN instrMgmt_dataOut[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.850 0.000 2004.130 4.000 ;
    END
  END instrMgmt_dataOut[19]
  PIN instrMgmt_dataOut[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.210 0.000 1896.490 4.000 ;
    END
  END instrMgmt_dataOut[1]
  PIN instrMgmt_dataOut[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.830 0.000 2010.110 4.000 ;
    END
  END instrMgmt_dataOut[20]
  PIN instrMgmt_dataOut[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END instrMgmt_dataOut[21]
  PIN instrMgmt_dataOut[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.790 0.000 2022.070 4.000 ;
    END
  END instrMgmt_dataOut[22]
  PIN instrMgmt_dataOut[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.770 0.000 2028.050 4.000 ;
    END
  END instrMgmt_dataOut[23]
  PIN instrMgmt_dataOut[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.750 0.000 2034.030 4.000 ;
    END
  END instrMgmt_dataOut[24]
  PIN instrMgmt_dataOut[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.730 0.000 2040.010 4.000 ;
    END
  END instrMgmt_dataOut[25]
  PIN instrMgmt_dataOut[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2045.710 0.000 2045.990 4.000 ;
    END
  END instrMgmt_dataOut[26]
  PIN instrMgmt_dataOut[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.690 0.000 2051.970 4.000 ;
    END
  END instrMgmt_dataOut[27]
  PIN instrMgmt_dataOut[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 0.000 2057.950 4.000 ;
    END
  END instrMgmt_dataOut[28]
  PIN instrMgmt_dataOut[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.650 0.000 2063.930 4.000 ;
    END
  END instrMgmt_dataOut[29]
  PIN instrMgmt_dataOut[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.190 0.000 1902.470 4.000 ;
    END
  END instrMgmt_dataOut[2]
  PIN instrMgmt_dataOut[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END instrMgmt_dataOut[30]
  PIN instrMgmt_dataOut[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.610 0.000 2075.890 4.000 ;
    END
  END instrMgmt_dataOut[31]
  PIN instrMgmt_dataOut[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.590 0.000 2081.870 4.000 ;
    END
  END instrMgmt_dataOut[32]
  PIN instrMgmt_dataOut[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2087.570 0.000 2087.850 4.000 ;
    END
  END instrMgmt_dataOut[33]
  PIN instrMgmt_dataOut[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.550 0.000 2093.830 4.000 ;
    END
  END instrMgmt_dataOut[34]
  PIN instrMgmt_dataOut[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 0.000 2099.810 4.000 ;
    END
  END instrMgmt_dataOut[35]
  PIN instrMgmt_dataOut[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.510 0.000 2105.790 4.000 ;
    END
  END instrMgmt_dataOut[36]
  PIN instrMgmt_dataOut[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.490 0.000 2111.770 4.000 ;
    END
  END instrMgmt_dataOut[37]
  PIN instrMgmt_dataOut[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.470 0.000 2117.750 4.000 ;
    END
  END instrMgmt_dataOut[38]
  PIN instrMgmt_dataOut[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2123.450 0.000 2123.730 4.000 ;
    END
  END instrMgmt_dataOut[39]
  PIN instrMgmt_dataOut[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.170 0.000 1908.450 4.000 ;
    END
  END instrMgmt_dataOut[3]
  PIN instrMgmt_dataOut[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.430 0.000 2129.710 4.000 ;
    END
  END instrMgmt_dataOut[40]
  PIN instrMgmt_dataOut[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.410 0.000 2135.690 4.000 ;
    END
  END instrMgmt_dataOut[41]
  PIN instrMgmt_dataOut[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END instrMgmt_dataOut[42]
  PIN instrMgmt_dataOut[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.370 0.000 2147.650 4.000 ;
    END
  END instrMgmt_dataOut[43]
  PIN instrMgmt_dataOut[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.350 0.000 2153.630 4.000 ;
    END
  END instrMgmt_dataOut[44]
  PIN instrMgmt_dataOut[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.330 0.000 2159.610 4.000 ;
    END
  END instrMgmt_dataOut[45]
  PIN instrMgmt_dataOut[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.310 0.000 2165.590 4.000 ;
    END
  END instrMgmt_dataOut[46]
  PIN instrMgmt_dataOut[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.290 0.000 2171.570 4.000 ;
    END
  END instrMgmt_dataOut[47]
  PIN instrMgmt_dataOut[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.270 0.000 2177.550 4.000 ;
    END
  END instrMgmt_dataOut[48]
  PIN instrMgmt_dataOut[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 0.000 2183.530 4.000 ;
    END
  END instrMgmt_dataOut[49]
  PIN instrMgmt_dataOut[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.150 0.000 1914.430 4.000 ;
    END
  END instrMgmt_dataOut[4]
  PIN instrMgmt_dataOut[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.230 0.000 2189.510 4.000 ;
    END
  END instrMgmt_dataOut[50]
  PIN instrMgmt_dataOut[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.210 0.000 2195.490 4.000 ;
    END
  END instrMgmt_dataOut[51]
  PIN instrMgmt_dataOut[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.190 0.000 2201.470 4.000 ;
    END
  END instrMgmt_dataOut[52]
  PIN instrMgmt_dataOut[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.170 0.000 2207.450 4.000 ;
    END
  END instrMgmt_dataOut[53]
  PIN instrMgmt_dataOut[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.150 0.000 2213.430 4.000 ;
    END
  END instrMgmt_dataOut[54]
  PIN instrMgmt_dataOut[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.130 0.000 2219.410 4.000 ;
    END
  END instrMgmt_dataOut[55]
  PIN instrMgmt_dataOut[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 0.000 2225.390 4.000 ;
    END
  END instrMgmt_dataOut[56]
  PIN instrMgmt_dataOut[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.090 0.000 2231.370 4.000 ;
    END
  END instrMgmt_dataOut[57]
  PIN instrMgmt_dataOut[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.070 0.000 2237.350 4.000 ;
    END
  END instrMgmt_dataOut[58]
  PIN instrMgmt_dataOut[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.050 0.000 2243.330 4.000 ;
    END
  END instrMgmt_dataOut[59]
  PIN instrMgmt_dataOut[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.130 0.000 1920.410 4.000 ;
    END
  END instrMgmt_dataOut[5]
  PIN instrMgmt_dataOut[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2249.030 0.000 2249.310 4.000 ;
    END
  END instrMgmt_dataOut[60]
  PIN instrMgmt_dataOut[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.010 0.000 2255.290 4.000 ;
    END
  END instrMgmt_dataOut[61]
  PIN instrMgmt_dataOut[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.990 0.000 2261.270 4.000 ;
    END
  END instrMgmt_dataOut[62]
  PIN instrMgmt_dataOut[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.970 0.000 2267.250 4.000 ;
    END
  END instrMgmt_dataOut[63]
  PIN instrMgmt_dataOut[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.110 0.000 1926.390 4.000 ;
    END
  END instrMgmt_dataOut[6]
  PIN instrMgmt_dataOut[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END instrMgmt_dataOut[7]
  PIN instrMgmt_dataOut[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 0.000 1938.350 4.000 ;
    END
  END instrMgmt_dataOut[8]
  PIN instrMgmt_dataOut[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.050 0.000 1944.330 4.000 ;
    END
  END instrMgmt_dataOut[9]
  PIN instrMgmt_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.930 0.000 2279.210 4.000 ;
    END
  END instrMgmt_we
  PIN instrMgmt_wm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.910 0.000 2285.190 4.000 ;
    END
  END instrMgmt_wm[0]
  PIN instrMgmt_wm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.890 0.000 2291.170 4.000 ;
    END
  END instrMgmt_wm[1]
  PIN instrMgmt_wm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2296.870 0.000 2297.150 4.000 ;
    END
  END instrMgmt_wm[2]
  PIN instrMgmt_wm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.850 0.000 2303.130 4.000 ;
    END
  END instrMgmt_wm[3]
  PIN instrMgmt_wm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.830 0.000 2309.110 4.000 ;
    END
  END instrMgmt_wm[4]
  PIN instrMgmt_wm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2314.810 0.000 2315.090 4.000 ;
    END
  END instrMgmt_wm[5]
  PIN instrMgmt_wm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.790 0.000 2321.070 4.000 ;
    END
  END instrMgmt_wm[6]
  PIN instrMgmt_wm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2326.770 0.000 2327.050 4.000 ;
    END
  END instrMgmt_wm[7]
  PIN instr_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.750 0.000 2333.030 4.000 ;
    END
  END instr_addr[0]
  PIN instr_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.730 0.000 2339.010 4.000 ;
    END
  END instr_addr[1]
  PIN instr_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.710 0.000 2344.990 4.000 ;
    END
  END instr_addr[2]
  PIN instr_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 0.000 2350.970 4.000 ;
    END
  END instr_addr[3]
  PIN instr_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.670 0.000 2356.950 4.000 ;
    END
  END instr_addr[4]
  PIN instr_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.650 0.000 2362.930 4.000 ;
    END
  END instr_addr[5]
  PIN instr_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.630 0.000 2368.910 4.000 ;
    END
  END instr_addr[6]
  PIN instr_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.610 0.000 2374.890 4.000 ;
    END
  END instr_addr[7]
  PIN instr_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2380.590 0.000 2380.870 4.000 ;
    END
  END instr_addr[8]
  PIN instr_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.290 0.000 2769.570 4.000 ;
    END
  END instr_ce
  PIN instr_dataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.570 0.000 2386.850 4.000 ;
    END
  END instr_dataIn[0]
  PIN instr_dataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.370 0.000 2446.650 4.000 ;
    END
  END instr_dataIn[10]
  PIN instr_dataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.350 0.000 2452.630 4.000 ;
    END
  END instr_dataIn[11]
  PIN instr_dataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.330 0.000 2458.610 4.000 ;
    END
  END instr_dataIn[12]
  PIN instr_dataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.310 0.000 2464.590 4.000 ;
    END
  END instr_dataIn[13]
  PIN instr_dataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.290 0.000 2470.570 4.000 ;
    END
  END instr_dataIn[14]
  PIN instr_dataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.270 0.000 2476.550 4.000 ;
    END
  END instr_dataIn[15]
  PIN instr_dataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.250 0.000 2482.530 4.000 ;
    END
  END instr_dataIn[16]
  PIN instr_dataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.230 0.000 2488.510 4.000 ;
    END
  END instr_dataIn[17]
  PIN instr_dataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.210 0.000 2494.490 4.000 ;
    END
  END instr_dataIn[18]
  PIN instr_dataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.190 0.000 2500.470 4.000 ;
    END
  END instr_dataIn[19]
  PIN instr_dataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 0.000 2392.830 4.000 ;
    END
  END instr_dataIn[1]
  PIN instr_dataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.170 0.000 2506.450 4.000 ;
    END
  END instr_dataIn[20]
  PIN instr_dataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.150 0.000 2512.430 4.000 ;
    END
  END instr_dataIn[21]
  PIN instr_dataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 0.000 2518.410 4.000 ;
    END
  END instr_dataIn[22]
  PIN instr_dataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2524.110 0.000 2524.390 4.000 ;
    END
  END instr_dataIn[23]
  PIN instr_dataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2530.090 0.000 2530.370 4.000 ;
    END
  END instr_dataIn[24]
  PIN instr_dataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2536.070 0.000 2536.350 4.000 ;
    END
  END instr_dataIn[25]
  PIN instr_dataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2542.050 0.000 2542.330 4.000 ;
    END
  END instr_dataIn[26]
  PIN instr_dataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2548.030 0.000 2548.310 4.000 ;
    END
  END instr_dataIn[27]
  PIN instr_dataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.010 0.000 2554.290 4.000 ;
    END
  END instr_dataIn[28]
  PIN instr_dataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.990 0.000 2560.270 4.000 ;
    END
  END instr_dataIn[29]
  PIN instr_dataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.530 0.000 2398.810 4.000 ;
    END
  END instr_dataIn[2]
  PIN instr_dataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.970 0.000 2566.250 4.000 ;
    END
  END instr_dataIn[30]
  PIN instr_dataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.950 0.000 2572.230 4.000 ;
    END
  END instr_dataIn[31]
  PIN instr_dataIn[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.930 0.000 2578.210 4.000 ;
    END
  END instr_dataIn[32]
  PIN instr_dataIn[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.910 0.000 2584.190 4.000 ;
    END
  END instr_dataIn[33]
  PIN instr_dataIn[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.890 0.000 2590.170 4.000 ;
    END
  END instr_dataIn[34]
  PIN instr_dataIn[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.870 0.000 2596.150 4.000 ;
    END
  END instr_dataIn[35]
  PIN instr_dataIn[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.850 0.000 2602.130 4.000 ;
    END
  END instr_dataIn[36]
  PIN instr_dataIn[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.830 0.000 2608.110 4.000 ;
    END
  END instr_dataIn[37]
  PIN instr_dataIn[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.810 0.000 2614.090 4.000 ;
    END
  END instr_dataIn[38]
  PIN instr_dataIn[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.790 0.000 2620.070 4.000 ;
    END
  END instr_dataIn[39]
  PIN instr_dataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2404.510 0.000 2404.790 4.000 ;
    END
  END instr_dataIn[3]
  PIN instr_dataIn[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.770 0.000 2626.050 4.000 ;
    END
  END instr_dataIn[40]
  PIN instr_dataIn[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.750 0.000 2632.030 4.000 ;
    END
  END instr_dataIn[41]
  PIN instr_dataIn[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.730 0.000 2638.010 4.000 ;
    END
  END instr_dataIn[42]
  PIN instr_dataIn[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.710 0.000 2643.990 4.000 ;
    END
  END instr_dataIn[43]
  PIN instr_dataIn[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.690 0.000 2649.970 4.000 ;
    END
  END instr_dataIn[44]
  PIN instr_dataIn[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.670 0.000 2655.950 4.000 ;
    END
  END instr_dataIn[45]
  PIN instr_dataIn[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.650 0.000 2661.930 4.000 ;
    END
  END instr_dataIn[46]
  PIN instr_dataIn[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.630 0.000 2667.910 4.000 ;
    END
  END instr_dataIn[47]
  PIN instr_dataIn[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2673.610 0.000 2673.890 4.000 ;
    END
  END instr_dataIn[48]
  PIN instr_dataIn[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2679.590 0.000 2679.870 4.000 ;
    END
  END instr_dataIn[49]
  PIN instr_dataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.490 0.000 2410.770 4.000 ;
    END
  END instr_dataIn[4]
  PIN instr_dataIn[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.570 0.000 2685.850 4.000 ;
    END
  END instr_dataIn[50]
  PIN instr_dataIn[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.550 0.000 2691.830 4.000 ;
    END
  END instr_dataIn[51]
  PIN instr_dataIn[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.530 0.000 2697.810 4.000 ;
    END
  END instr_dataIn[52]
  PIN instr_dataIn[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.510 0.000 2703.790 4.000 ;
    END
  END instr_dataIn[53]
  PIN instr_dataIn[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.490 0.000 2709.770 4.000 ;
    END
  END instr_dataIn[54]
  PIN instr_dataIn[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.470 0.000 2715.750 4.000 ;
    END
  END instr_dataIn[55]
  PIN instr_dataIn[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.450 0.000 2721.730 4.000 ;
    END
  END instr_dataIn[56]
  PIN instr_dataIn[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.430 0.000 2727.710 4.000 ;
    END
  END instr_dataIn[57]
  PIN instr_dataIn[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.410 0.000 2733.690 4.000 ;
    END
  END instr_dataIn[58]
  PIN instr_dataIn[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.390 0.000 2739.670 4.000 ;
    END
  END instr_dataIn[59]
  PIN instr_dataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.470 0.000 2416.750 4.000 ;
    END
  END instr_dataIn[5]
  PIN instr_dataIn[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.370 0.000 2745.650 4.000 ;
    END
  END instr_dataIn[60]
  PIN instr_dataIn[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.350 0.000 2751.630 4.000 ;
    END
  END instr_dataIn[61]
  PIN instr_dataIn[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.330 0.000 2757.610 4.000 ;
    END
  END instr_dataIn[62]
  PIN instr_dataIn[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.310 0.000 2763.590 4.000 ;
    END
  END instr_dataIn[63]
  PIN instr_dataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.450 0.000 2422.730 4.000 ;
    END
  END instr_dataIn[6]
  PIN instr_dataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.430 0.000 2428.710 4.000 ;
    END
  END instr_dataIn[7]
  PIN instr_dataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 0.000 2434.690 4.000 ;
    END
  END instr_dataIn[8]
  PIN instr_dataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.390 0.000 2440.670 4.000 ;
    END
  END instr_dataIn[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 29.280 2800.000 29.880 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1436.880 2800.000 1437.480 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1577.640 2800.000 1578.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1718.400 2800.000 1719.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1859.160 2800.000 1859.760 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1999.920 2800.000 2000.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.350 2496.000 2153.630 2500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 2496.000 2225.390 2500.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2296.870 2496.000 2297.150 2500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.630 2496.000 2368.910 2500.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.390 2496.000 2440.670 2500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 170.040 2800.000 170.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.150 2496.000 2512.430 2500.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.910 2496.000 2584.190 2500.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.670 2496.000 2655.950 2500.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.430 2496.000 2727.710 2500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 310.800 2800.000 311.400 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1133.600 4.000 1134.200 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1549.760 4.000 1550.360 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1688.480 4.000 1689.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1827.200 4.000 1827.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 451.560 2800.000 452.160 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 592.320 2800.000 592.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 733.080 2800.000 733.680 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 873.840 2800.000 874.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1014.600 2800.000 1015.200 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1155.360 2800.000 1155.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1296.120 2800.000 1296.720 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 76.200 2800.000 76.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1483.800 2800.000 1484.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1624.560 2800.000 1625.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1765.320 2800.000 1765.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1906.080 2800.000 1906.680 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2046.840 2800.000 2047.440 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.270 2496.000 2177.550 2500.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2249.030 2496.000 2249.310 2500.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.790 2496.000 2321.070 2500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 2496.000 2392.830 2500.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.310 2496.000 2464.590 2500.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 216.960 2800.000 217.560 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2536.070 2496.000 2536.350 2500.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.830 2496.000 2608.110 2500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2679.590 2496.000 2679.870 2500.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.350 2496.000 2751.630 2500.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.680 4.000 764.280 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 357.720 2800.000 358.320 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1318.560 4.000 1319.160 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.280 4.000 1457.880 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.000 4.000 1596.600 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.720 4.000 1735.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1873.440 4.000 1874.040 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 498.480 2800.000 499.080 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 639.240 2800.000 639.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 780.000 2800.000 780.600 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 920.760 2800.000 921.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1061.520 2800.000 1062.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1202.280 2800.000 1202.880 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1343.040 2800.000 1343.640 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 123.120 2800.000 123.720 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1530.720 2800.000 1531.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1671.480 2800.000 1672.080 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1812.240 2800.000 1812.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1953.000 2800.000 1953.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 2093.760 2800.000 2094.360 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.190 2496.000 2201.470 2500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.950 2496.000 2273.230 2500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.710 2496.000 2344.990 2500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.470 2496.000 2416.750 2500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.230 2496.000 2488.510 2500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 263.880 2800.000 264.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.990 2496.000 2560.270 2500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.750 2496.000 2632.030 2500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.510 2496.000 2703.790 2500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2775.270 2496.000 2775.550 2500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 404.640 2800.000 405.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1226.080 4.000 1226.680 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.800 4.000 1365.400 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1503.520 4.000 1504.120 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1642.240 4.000 1642.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1780.960 4.000 1781.560 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1919.680 4.000 1920.280 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 545.400 2800.000 546.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 686.160 2800.000 686.760 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 826.920 2800.000 827.520 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 967.680 2800.000 968.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1108.440 2800.000 1109.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1249.200 2800.000 1249.800 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1389.960 2800.000 1390.560 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END irq[2]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 0.000 1286.530 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230 0.000 1292.510 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 0.000 1310.450 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 0.000 1322.410 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 0.000 1328.390 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 0.000 1334.370 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 0.000 1340.350 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.030 0.000 1352.310 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 0.000 1358.290 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.970 0.000 1370.250 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 0.000 1412.110 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 0.000 1424.070 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 0.000 1436.030 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 0.000 1442.010 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 0.000 873.910 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 0.000 975.570 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 0.000 981.550 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 0.000 1041.350 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 0.000 1101.150 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 0.000 1119.090 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 0.000 1143.010 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 0.000 1148.990 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 0.000 1166.930 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 0.000 1172.910 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.590 0.000 1184.870 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.570 0.000 1190.850 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 0.000 1196.830 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 0.000 1202.810 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 0.000 1214.770 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 0.000 1244.670 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 0.000 1268.590 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END la_data_out[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 2496.000 24.750 2500.000 ;
    END
  END mem_addr[0]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 2496.000 48.670 2500.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 2496.000 72.590 2500.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 2496.000 96.510 2500.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 2496.000 120.430 2500.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 2496.000 144.350 2500.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 2496.000 168.270 2500.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 2496.000 192.190 2500.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 2496.000 216.110 2500.000 ;
    END
  END mem_addr[8]
  PIN mem_ce
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 2496.000 1890.510 2500.000 ;
    END
  END mem_ce
  PIN mem_dataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 2496.000 240.030 2500.000 ;
    END
  END mem_dataIn[0]
  PIN mem_dataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 2496.000 479.230 2500.000 ;
    END
  END mem_dataIn[10]
  PIN mem_dataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 2496.000 503.150 2500.000 ;
    END
  END mem_dataIn[11]
  PIN mem_dataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 2496.000 527.070 2500.000 ;
    END
  END mem_dataIn[12]
  PIN mem_dataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 2496.000 550.990 2500.000 ;
    END
  END mem_dataIn[13]
  PIN mem_dataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 2496.000 574.910 2500.000 ;
    END
  END mem_dataIn[14]
  PIN mem_dataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 2496.000 598.830 2500.000 ;
    END
  END mem_dataIn[15]
  PIN mem_dataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 2496.000 622.750 2500.000 ;
    END
  END mem_dataIn[16]
  PIN mem_dataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 2496.000 646.670 2500.000 ;
    END
  END mem_dataIn[17]
  PIN mem_dataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 2496.000 670.590 2500.000 ;
    END
  END mem_dataIn[18]
  PIN mem_dataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 2496.000 694.510 2500.000 ;
    END
  END mem_dataIn[19]
  PIN mem_dataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 2496.000 263.950 2500.000 ;
    END
  END mem_dataIn[1]
  PIN mem_dataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 2496.000 718.430 2500.000 ;
    END
  END mem_dataIn[20]
  PIN mem_dataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 2496.000 742.350 2500.000 ;
    END
  END mem_dataIn[21]
  PIN mem_dataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 2496.000 766.270 2500.000 ;
    END
  END mem_dataIn[22]
  PIN mem_dataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 2496.000 790.190 2500.000 ;
    END
  END mem_dataIn[23]
  PIN mem_dataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 2496.000 814.110 2500.000 ;
    END
  END mem_dataIn[24]
  PIN mem_dataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 2496.000 838.030 2500.000 ;
    END
  END mem_dataIn[25]
  PIN mem_dataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 2496.000 861.950 2500.000 ;
    END
  END mem_dataIn[26]
  PIN mem_dataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 2496.000 885.870 2500.000 ;
    END
  END mem_dataIn[27]
  PIN mem_dataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 2496.000 909.790 2500.000 ;
    END
  END mem_dataIn[28]
  PIN mem_dataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 2496.000 933.710 2500.000 ;
    END
  END mem_dataIn[29]
  PIN mem_dataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 2496.000 287.870 2500.000 ;
    END
  END mem_dataIn[2]
  PIN mem_dataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 2496.000 957.630 2500.000 ;
    END
  END mem_dataIn[30]
  PIN mem_dataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 2496.000 981.550 2500.000 ;
    END
  END mem_dataIn[31]
  PIN mem_dataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 2496.000 311.790 2500.000 ;
    END
  END mem_dataIn[3]
  PIN mem_dataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 2496.000 335.710 2500.000 ;
    END
  END mem_dataIn[4]
  PIN mem_dataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 2496.000 359.630 2500.000 ;
    END
  END mem_dataIn[5]
  PIN mem_dataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 2496.000 383.550 2500.000 ;
    END
  END mem_dataIn[6]
  PIN mem_dataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 2496.000 407.470 2500.000 ;
    END
  END mem_dataIn[7]
  PIN mem_dataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 2496.000 431.390 2500.000 ;
    END
  END mem_dataIn[8]
  PIN mem_dataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 2496.000 455.310 2500.000 ;
    END
  END mem_dataIn[9]
  PIN mem_dataOut[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 2496.000 1005.470 2500.000 ;
    END
  END mem_dataOut[0]
  PIN mem_dataOut[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.390 2496.000 1244.670 2500.000 ;
    END
  END mem_dataOut[10]
  PIN mem_dataOut[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 2496.000 1268.590 2500.000 ;
    END
  END mem_dataOut[11]
  PIN mem_dataOut[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230 2496.000 1292.510 2500.000 ;
    END
  END mem_dataOut[12]
  PIN mem_dataOut[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 2496.000 1316.430 2500.000 ;
    END
  END mem_dataOut[13]
  PIN mem_dataOut[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 2496.000 1340.350 2500.000 ;
    END
  END mem_dataOut[14]
  PIN mem_dataOut[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 2496.000 1364.270 2500.000 ;
    END
  END mem_dataOut[15]
  PIN mem_dataOut[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 2496.000 1388.190 2500.000 ;
    END
  END mem_dataOut[16]
  PIN mem_dataOut[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 2496.000 1412.110 2500.000 ;
    END
  END mem_dataOut[17]
  PIN mem_dataOut[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 2496.000 1436.030 2500.000 ;
    END
  END mem_dataOut[18]
  PIN mem_dataOut[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 2496.000 1459.950 2500.000 ;
    END
  END mem_dataOut[19]
  PIN mem_dataOut[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 2496.000 1029.390 2500.000 ;
    END
  END mem_dataOut[1]
  PIN mem_dataOut[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 2496.000 1483.870 2500.000 ;
    END
  END mem_dataOut[20]
  PIN mem_dataOut[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 2496.000 1507.790 2500.000 ;
    END
  END mem_dataOut[21]
  PIN mem_dataOut[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.430 2496.000 1531.710 2500.000 ;
    END
  END mem_dataOut[22]
  PIN mem_dataOut[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 2496.000 1555.630 2500.000 ;
    END
  END mem_dataOut[23]
  PIN mem_dataOut[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 2496.000 1579.550 2500.000 ;
    END
  END mem_dataOut[24]
  PIN mem_dataOut[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.190 2496.000 1603.470 2500.000 ;
    END
  END mem_dataOut[25]
  PIN mem_dataOut[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 2496.000 1627.390 2500.000 ;
    END
  END mem_dataOut[26]
  PIN mem_dataOut[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 2496.000 1651.310 2500.000 ;
    END
  END mem_dataOut[27]
  PIN mem_dataOut[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 2496.000 1675.230 2500.000 ;
    END
  END mem_dataOut[28]
  PIN mem_dataOut[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 2496.000 1699.150 2500.000 ;
    END
  END mem_dataOut[29]
  PIN mem_dataOut[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 2496.000 1053.310 2500.000 ;
    END
  END mem_dataOut[2]
  PIN mem_dataOut[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 2496.000 1723.070 2500.000 ;
    END
  END mem_dataOut[30]
  PIN mem_dataOut[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.710 2496.000 1746.990 2500.000 ;
    END
  END mem_dataOut[31]
  PIN mem_dataOut[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 2496.000 1077.230 2500.000 ;
    END
  END mem_dataOut[3]
  PIN mem_dataOut[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 2496.000 1101.150 2500.000 ;
    END
  END mem_dataOut[4]
  PIN mem_dataOut[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 2496.000 1125.070 2500.000 ;
    END
  END mem_dataOut[5]
  PIN mem_dataOut[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 2496.000 1148.990 2500.000 ;
    END
  END mem_dataOut[6]
  PIN mem_dataOut[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 2496.000 1172.910 2500.000 ;
    END
  END mem_dataOut[7]
  PIN mem_dataOut[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.550 2496.000 1196.830 2500.000 ;
    END
  END mem_dataOut[8]
  PIN mem_dataOut[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 2496.000 1220.750 2500.000 ;
    END
  END mem_dataOut[9]
  PIN mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.310 2496.000 1866.590 2500.000 ;
    END
  END mem_we
  PIN mem_wm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 2496.000 1770.910 2500.000 ;
    END
  END mem_wm[0]
  PIN mem_wm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.550 2496.000 1794.830 2500.000 ;
    END
  END mem_wm[1]
  PIN mem_wm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.470 2496.000 1818.750 2500.000 ;
    END
  END mem_wm[2]
  PIN mem_wm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.390 2496.000 1842.670 2500.000 ;
    END
  END mem_wm[3]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 2489.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 2489.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.150 2496.000 1914.430 2500.000 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 2488.885 ;
      LAYER met1 ;
        RECT 5.520 0.720 2794.040 2497.940 ;
      LAYER met2 ;
        RECT 7.910 2495.720 24.190 2497.970 ;
        RECT 25.030 2495.720 48.110 2497.970 ;
        RECT 48.950 2495.720 72.030 2497.970 ;
        RECT 72.870 2495.720 95.950 2497.970 ;
        RECT 96.790 2495.720 119.870 2497.970 ;
        RECT 120.710 2495.720 143.790 2497.970 ;
        RECT 144.630 2495.720 167.710 2497.970 ;
        RECT 168.550 2495.720 191.630 2497.970 ;
        RECT 192.470 2495.720 215.550 2497.970 ;
        RECT 216.390 2495.720 239.470 2497.970 ;
        RECT 240.310 2495.720 263.390 2497.970 ;
        RECT 264.230 2495.720 287.310 2497.970 ;
        RECT 288.150 2495.720 311.230 2497.970 ;
        RECT 312.070 2495.720 335.150 2497.970 ;
        RECT 335.990 2495.720 359.070 2497.970 ;
        RECT 359.910 2495.720 382.990 2497.970 ;
        RECT 383.830 2495.720 406.910 2497.970 ;
        RECT 407.750 2495.720 430.830 2497.970 ;
        RECT 431.670 2495.720 454.750 2497.970 ;
        RECT 455.590 2495.720 478.670 2497.970 ;
        RECT 479.510 2495.720 502.590 2497.970 ;
        RECT 503.430 2495.720 526.510 2497.970 ;
        RECT 527.350 2495.720 550.430 2497.970 ;
        RECT 551.270 2495.720 574.350 2497.970 ;
        RECT 575.190 2495.720 598.270 2497.970 ;
        RECT 599.110 2495.720 622.190 2497.970 ;
        RECT 623.030 2495.720 646.110 2497.970 ;
        RECT 646.950 2495.720 670.030 2497.970 ;
        RECT 670.870 2495.720 693.950 2497.970 ;
        RECT 694.790 2495.720 717.870 2497.970 ;
        RECT 718.710 2495.720 741.790 2497.970 ;
        RECT 742.630 2495.720 765.710 2497.970 ;
        RECT 766.550 2495.720 789.630 2497.970 ;
        RECT 790.470 2495.720 813.550 2497.970 ;
        RECT 814.390 2495.720 837.470 2497.970 ;
        RECT 838.310 2495.720 861.390 2497.970 ;
        RECT 862.230 2495.720 885.310 2497.970 ;
        RECT 886.150 2495.720 909.230 2497.970 ;
        RECT 910.070 2495.720 933.150 2497.970 ;
        RECT 933.990 2495.720 957.070 2497.970 ;
        RECT 957.910 2495.720 980.990 2497.970 ;
        RECT 981.830 2495.720 1004.910 2497.970 ;
        RECT 1005.750 2495.720 1028.830 2497.970 ;
        RECT 1029.670 2495.720 1052.750 2497.970 ;
        RECT 1053.590 2495.720 1076.670 2497.970 ;
        RECT 1077.510 2495.720 1100.590 2497.970 ;
        RECT 1101.430 2495.720 1124.510 2497.970 ;
        RECT 1125.350 2495.720 1148.430 2497.970 ;
        RECT 1149.270 2495.720 1172.350 2497.970 ;
        RECT 1173.190 2495.720 1196.270 2497.970 ;
        RECT 1197.110 2495.720 1220.190 2497.970 ;
        RECT 1221.030 2495.720 1244.110 2497.970 ;
        RECT 1244.950 2495.720 1268.030 2497.970 ;
        RECT 1268.870 2495.720 1291.950 2497.970 ;
        RECT 1292.790 2495.720 1315.870 2497.970 ;
        RECT 1316.710 2495.720 1339.790 2497.970 ;
        RECT 1340.630 2495.720 1363.710 2497.970 ;
        RECT 1364.550 2495.720 1387.630 2497.970 ;
        RECT 1388.470 2495.720 1411.550 2497.970 ;
        RECT 1412.390 2495.720 1435.470 2497.970 ;
        RECT 1436.310 2495.720 1459.390 2497.970 ;
        RECT 1460.230 2495.720 1483.310 2497.970 ;
        RECT 1484.150 2495.720 1507.230 2497.970 ;
        RECT 1508.070 2495.720 1531.150 2497.970 ;
        RECT 1531.990 2495.720 1555.070 2497.970 ;
        RECT 1555.910 2495.720 1578.990 2497.970 ;
        RECT 1579.830 2495.720 1602.910 2497.970 ;
        RECT 1603.750 2495.720 1626.830 2497.970 ;
        RECT 1627.670 2495.720 1650.750 2497.970 ;
        RECT 1651.590 2495.720 1674.670 2497.970 ;
        RECT 1675.510 2495.720 1698.590 2497.970 ;
        RECT 1699.430 2495.720 1722.510 2497.970 ;
        RECT 1723.350 2495.720 1746.430 2497.970 ;
        RECT 1747.270 2495.720 1770.350 2497.970 ;
        RECT 1771.190 2495.720 1794.270 2497.970 ;
        RECT 1795.110 2495.720 1818.190 2497.970 ;
        RECT 1819.030 2495.720 1842.110 2497.970 ;
        RECT 1842.950 2495.720 1866.030 2497.970 ;
        RECT 1866.870 2495.720 1889.950 2497.970 ;
        RECT 1890.790 2495.720 1913.870 2497.970 ;
        RECT 1914.710 2495.720 1937.790 2497.970 ;
        RECT 1938.630 2495.720 1961.710 2497.970 ;
        RECT 1962.550 2495.720 1985.630 2497.970 ;
        RECT 1986.470 2495.720 2009.550 2497.970 ;
        RECT 2010.390 2495.720 2033.470 2497.970 ;
        RECT 2034.310 2495.720 2057.390 2497.970 ;
        RECT 2058.230 2495.720 2081.310 2497.970 ;
        RECT 2082.150 2495.720 2105.230 2497.970 ;
        RECT 2106.070 2495.720 2129.150 2497.970 ;
        RECT 2129.990 2495.720 2153.070 2497.970 ;
        RECT 2153.910 2495.720 2176.990 2497.970 ;
        RECT 2177.830 2495.720 2200.910 2497.970 ;
        RECT 2201.750 2495.720 2224.830 2497.970 ;
        RECT 2225.670 2495.720 2248.750 2497.970 ;
        RECT 2249.590 2495.720 2272.670 2497.970 ;
        RECT 2273.510 2495.720 2296.590 2497.970 ;
        RECT 2297.430 2495.720 2320.510 2497.970 ;
        RECT 2321.350 2495.720 2344.430 2497.970 ;
        RECT 2345.270 2495.720 2368.350 2497.970 ;
        RECT 2369.190 2495.720 2392.270 2497.970 ;
        RECT 2393.110 2495.720 2416.190 2497.970 ;
        RECT 2417.030 2495.720 2440.110 2497.970 ;
        RECT 2440.950 2495.720 2464.030 2497.970 ;
        RECT 2464.870 2495.720 2487.950 2497.970 ;
        RECT 2488.790 2495.720 2511.870 2497.970 ;
        RECT 2512.710 2495.720 2535.790 2497.970 ;
        RECT 2536.630 2495.720 2559.710 2497.970 ;
        RECT 2560.550 2495.720 2583.630 2497.970 ;
        RECT 2584.470 2495.720 2607.550 2497.970 ;
        RECT 2608.390 2495.720 2631.470 2497.970 ;
        RECT 2632.310 2495.720 2655.390 2497.970 ;
        RECT 2656.230 2495.720 2679.310 2497.970 ;
        RECT 2680.150 2495.720 2703.230 2497.970 ;
        RECT 2704.070 2495.720 2727.150 2497.970 ;
        RECT 2727.990 2495.720 2751.070 2497.970 ;
        RECT 2751.910 2495.720 2774.990 2497.970 ;
        RECT 2775.830 2495.720 2792.560 2497.970 ;
        RECT 7.910 4.280 2792.560 2495.720 ;
        RECT 7.910 0.690 30.170 4.280 ;
        RECT 31.010 0.690 36.150 4.280 ;
        RECT 36.990 0.690 42.130 4.280 ;
        RECT 42.970 0.690 48.110 4.280 ;
        RECT 48.950 0.690 54.090 4.280 ;
        RECT 54.930 0.690 60.070 4.280 ;
        RECT 60.910 0.690 66.050 4.280 ;
        RECT 66.890 0.690 72.030 4.280 ;
        RECT 72.870 0.690 78.010 4.280 ;
        RECT 78.850 0.690 83.990 4.280 ;
        RECT 84.830 0.690 89.970 4.280 ;
        RECT 90.810 0.690 95.950 4.280 ;
        RECT 96.790 0.690 101.930 4.280 ;
        RECT 102.770 0.690 107.910 4.280 ;
        RECT 108.750 0.690 113.890 4.280 ;
        RECT 114.730 0.690 119.870 4.280 ;
        RECT 120.710 0.690 125.850 4.280 ;
        RECT 126.690 0.690 131.830 4.280 ;
        RECT 132.670 0.690 137.810 4.280 ;
        RECT 138.650 0.690 143.790 4.280 ;
        RECT 144.630 0.690 149.770 4.280 ;
        RECT 150.610 0.690 155.750 4.280 ;
        RECT 156.590 0.690 161.730 4.280 ;
        RECT 162.570 0.690 167.710 4.280 ;
        RECT 168.550 0.690 173.690 4.280 ;
        RECT 174.530 0.690 179.670 4.280 ;
        RECT 180.510 0.690 185.650 4.280 ;
        RECT 186.490 0.690 191.630 4.280 ;
        RECT 192.470 0.690 197.610 4.280 ;
        RECT 198.450 0.690 203.590 4.280 ;
        RECT 204.430 0.690 209.570 4.280 ;
        RECT 210.410 0.690 215.550 4.280 ;
        RECT 216.390 0.690 221.530 4.280 ;
        RECT 222.370 0.690 227.510 4.280 ;
        RECT 228.350 0.690 233.490 4.280 ;
        RECT 234.330 0.690 239.470 4.280 ;
        RECT 240.310 0.690 245.450 4.280 ;
        RECT 246.290 0.690 251.430 4.280 ;
        RECT 252.270 0.690 257.410 4.280 ;
        RECT 258.250 0.690 263.390 4.280 ;
        RECT 264.230 0.690 269.370 4.280 ;
        RECT 270.210 0.690 275.350 4.280 ;
        RECT 276.190 0.690 281.330 4.280 ;
        RECT 282.170 0.690 287.310 4.280 ;
        RECT 288.150 0.690 293.290 4.280 ;
        RECT 294.130 0.690 299.270 4.280 ;
        RECT 300.110 0.690 305.250 4.280 ;
        RECT 306.090 0.690 311.230 4.280 ;
        RECT 312.070 0.690 317.210 4.280 ;
        RECT 318.050 0.690 323.190 4.280 ;
        RECT 324.030 0.690 329.170 4.280 ;
        RECT 330.010 0.690 335.150 4.280 ;
        RECT 335.990 0.690 341.130 4.280 ;
        RECT 341.970 0.690 347.110 4.280 ;
        RECT 347.950 0.690 353.090 4.280 ;
        RECT 353.930 0.690 359.070 4.280 ;
        RECT 359.910 0.690 365.050 4.280 ;
        RECT 365.890 0.690 371.030 4.280 ;
        RECT 371.870 0.690 377.010 4.280 ;
        RECT 377.850 0.690 382.990 4.280 ;
        RECT 383.830 0.690 388.970 4.280 ;
        RECT 389.810 0.690 394.950 4.280 ;
        RECT 395.790 0.690 400.930 4.280 ;
        RECT 401.770 0.690 406.910 4.280 ;
        RECT 407.750 0.690 412.890 4.280 ;
        RECT 413.730 0.690 418.870 4.280 ;
        RECT 419.710 0.690 424.850 4.280 ;
        RECT 425.690 0.690 430.830 4.280 ;
        RECT 431.670 0.690 436.810 4.280 ;
        RECT 437.650 0.690 442.790 4.280 ;
        RECT 443.630 0.690 448.770 4.280 ;
        RECT 449.610 0.690 454.750 4.280 ;
        RECT 455.590 0.690 460.730 4.280 ;
        RECT 461.570 0.690 466.710 4.280 ;
        RECT 467.550 0.690 472.690 4.280 ;
        RECT 473.530 0.690 478.670 4.280 ;
        RECT 479.510 0.690 484.650 4.280 ;
        RECT 485.490 0.690 490.630 4.280 ;
        RECT 491.470 0.690 496.610 4.280 ;
        RECT 497.450 0.690 502.590 4.280 ;
        RECT 503.430 0.690 508.570 4.280 ;
        RECT 509.410 0.690 514.550 4.280 ;
        RECT 515.390 0.690 520.530 4.280 ;
        RECT 521.370 0.690 526.510 4.280 ;
        RECT 527.350 0.690 532.490 4.280 ;
        RECT 533.330 0.690 538.470 4.280 ;
        RECT 539.310 0.690 544.450 4.280 ;
        RECT 545.290 0.690 550.430 4.280 ;
        RECT 551.270 0.690 556.410 4.280 ;
        RECT 557.250 0.690 562.390 4.280 ;
        RECT 563.230 0.690 568.370 4.280 ;
        RECT 569.210 0.690 574.350 4.280 ;
        RECT 575.190 0.690 580.330 4.280 ;
        RECT 581.170 0.690 586.310 4.280 ;
        RECT 587.150 0.690 592.290 4.280 ;
        RECT 593.130 0.690 598.270 4.280 ;
        RECT 599.110 0.690 604.250 4.280 ;
        RECT 605.090 0.690 610.230 4.280 ;
        RECT 611.070 0.690 616.210 4.280 ;
        RECT 617.050 0.690 622.190 4.280 ;
        RECT 623.030 0.690 628.170 4.280 ;
        RECT 629.010 0.690 634.150 4.280 ;
        RECT 634.990 0.690 640.130 4.280 ;
        RECT 640.970 0.690 646.110 4.280 ;
        RECT 646.950 0.690 652.090 4.280 ;
        RECT 652.930 0.690 658.070 4.280 ;
        RECT 658.910 0.690 664.050 4.280 ;
        RECT 664.890 0.690 670.030 4.280 ;
        RECT 670.870 0.690 676.010 4.280 ;
        RECT 676.850 0.690 681.990 4.280 ;
        RECT 682.830 0.690 687.970 4.280 ;
        RECT 688.810 0.690 693.950 4.280 ;
        RECT 694.790 0.690 699.930 4.280 ;
        RECT 700.770 0.690 705.910 4.280 ;
        RECT 706.750 0.690 711.890 4.280 ;
        RECT 712.730 0.690 717.870 4.280 ;
        RECT 718.710 0.690 723.850 4.280 ;
        RECT 724.690 0.690 729.830 4.280 ;
        RECT 730.670 0.690 735.810 4.280 ;
        RECT 736.650 0.690 741.790 4.280 ;
        RECT 742.630 0.690 747.770 4.280 ;
        RECT 748.610 0.690 753.750 4.280 ;
        RECT 754.590 0.690 759.730 4.280 ;
        RECT 760.570 0.690 765.710 4.280 ;
        RECT 766.550 0.690 771.690 4.280 ;
        RECT 772.530 0.690 777.670 4.280 ;
        RECT 778.510 0.690 783.650 4.280 ;
        RECT 784.490 0.690 789.630 4.280 ;
        RECT 790.470 0.690 795.610 4.280 ;
        RECT 796.450 0.690 801.590 4.280 ;
        RECT 802.430 0.690 807.570 4.280 ;
        RECT 808.410 0.690 813.550 4.280 ;
        RECT 814.390 0.690 819.530 4.280 ;
        RECT 820.370 0.690 825.510 4.280 ;
        RECT 826.350 0.690 831.490 4.280 ;
        RECT 832.330 0.690 837.470 4.280 ;
        RECT 838.310 0.690 843.450 4.280 ;
        RECT 844.290 0.690 849.430 4.280 ;
        RECT 850.270 0.690 855.410 4.280 ;
        RECT 856.250 0.690 861.390 4.280 ;
        RECT 862.230 0.690 867.370 4.280 ;
        RECT 868.210 0.690 873.350 4.280 ;
        RECT 874.190 0.690 879.330 4.280 ;
        RECT 880.170 0.690 885.310 4.280 ;
        RECT 886.150 0.690 891.290 4.280 ;
        RECT 892.130 0.690 897.270 4.280 ;
        RECT 898.110 0.690 903.250 4.280 ;
        RECT 904.090 0.690 909.230 4.280 ;
        RECT 910.070 0.690 915.210 4.280 ;
        RECT 916.050 0.690 921.190 4.280 ;
        RECT 922.030 0.690 927.170 4.280 ;
        RECT 928.010 0.690 933.150 4.280 ;
        RECT 933.990 0.690 939.130 4.280 ;
        RECT 939.970 0.690 945.110 4.280 ;
        RECT 945.950 0.690 951.090 4.280 ;
        RECT 951.930 0.690 957.070 4.280 ;
        RECT 957.910 0.690 963.050 4.280 ;
        RECT 963.890 0.690 969.030 4.280 ;
        RECT 969.870 0.690 975.010 4.280 ;
        RECT 975.850 0.690 980.990 4.280 ;
        RECT 981.830 0.690 986.970 4.280 ;
        RECT 987.810 0.690 992.950 4.280 ;
        RECT 993.790 0.690 998.930 4.280 ;
        RECT 999.770 0.690 1004.910 4.280 ;
        RECT 1005.750 0.690 1010.890 4.280 ;
        RECT 1011.730 0.690 1016.870 4.280 ;
        RECT 1017.710 0.690 1022.850 4.280 ;
        RECT 1023.690 0.690 1028.830 4.280 ;
        RECT 1029.670 0.690 1034.810 4.280 ;
        RECT 1035.650 0.690 1040.790 4.280 ;
        RECT 1041.630 0.690 1046.770 4.280 ;
        RECT 1047.610 0.690 1052.750 4.280 ;
        RECT 1053.590 0.690 1058.730 4.280 ;
        RECT 1059.570 0.690 1064.710 4.280 ;
        RECT 1065.550 0.690 1070.690 4.280 ;
        RECT 1071.530 0.690 1076.670 4.280 ;
        RECT 1077.510 0.690 1082.650 4.280 ;
        RECT 1083.490 0.690 1088.630 4.280 ;
        RECT 1089.470 0.690 1094.610 4.280 ;
        RECT 1095.450 0.690 1100.590 4.280 ;
        RECT 1101.430 0.690 1106.570 4.280 ;
        RECT 1107.410 0.690 1112.550 4.280 ;
        RECT 1113.390 0.690 1118.530 4.280 ;
        RECT 1119.370 0.690 1124.510 4.280 ;
        RECT 1125.350 0.690 1130.490 4.280 ;
        RECT 1131.330 0.690 1136.470 4.280 ;
        RECT 1137.310 0.690 1142.450 4.280 ;
        RECT 1143.290 0.690 1148.430 4.280 ;
        RECT 1149.270 0.690 1154.410 4.280 ;
        RECT 1155.250 0.690 1160.390 4.280 ;
        RECT 1161.230 0.690 1166.370 4.280 ;
        RECT 1167.210 0.690 1172.350 4.280 ;
        RECT 1173.190 0.690 1178.330 4.280 ;
        RECT 1179.170 0.690 1184.310 4.280 ;
        RECT 1185.150 0.690 1190.290 4.280 ;
        RECT 1191.130 0.690 1196.270 4.280 ;
        RECT 1197.110 0.690 1202.250 4.280 ;
        RECT 1203.090 0.690 1208.230 4.280 ;
        RECT 1209.070 0.690 1214.210 4.280 ;
        RECT 1215.050 0.690 1220.190 4.280 ;
        RECT 1221.030 0.690 1226.170 4.280 ;
        RECT 1227.010 0.690 1232.150 4.280 ;
        RECT 1232.990 0.690 1238.130 4.280 ;
        RECT 1238.970 0.690 1244.110 4.280 ;
        RECT 1244.950 0.690 1250.090 4.280 ;
        RECT 1250.930 0.690 1256.070 4.280 ;
        RECT 1256.910 0.690 1262.050 4.280 ;
        RECT 1262.890 0.690 1268.030 4.280 ;
        RECT 1268.870 0.690 1274.010 4.280 ;
        RECT 1274.850 0.690 1279.990 4.280 ;
        RECT 1280.830 0.690 1285.970 4.280 ;
        RECT 1286.810 0.690 1291.950 4.280 ;
        RECT 1292.790 0.690 1297.930 4.280 ;
        RECT 1298.770 0.690 1303.910 4.280 ;
        RECT 1304.750 0.690 1309.890 4.280 ;
        RECT 1310.730 0.690 1315.870 4.280 ;
        RECT 1316.710 0.690 1321.850 4.280 ;
        RECT 1322.690 0.690 1327.830 4.280 ;
        RECT 1328.670 0.690 1333.810 4.280 ;
        RECT 1334.650 0.690 1339.790 4.280 ;
        RECT 1340.630 0.690 1345.770 4.280 ;
        RECT 1346.610 0.690 1351.750 4.280 ;
        RECT 1352.590 0.690 1357.730 4.280 ;
        RECT 1358.570 0.690 1363.710 4.280 ;
        RECT 1364.550 0.690 1369.690 4.280 ;
        RECT 1370.530 0.690 1375.670 4.280 ;
        RECT 1376.510 0.690 1381.650 4.280 ;
        RECT 1382.490 0.690 1387.630 4.280 ;
        RECT 1388.470 0.690 1393.610 4.280 ;
        RECT 1394.450 0.690 1399.590 4.280 ;
        RECT 1400.430 0.690 1405.570 4.280 ;
        RECT 1406.410 0.690 1411.550 4.280 ;
        RECT 1412.390 0.690 1417.530 4.280 ;
        RECT 1418.370 0.690 1423.510 4.280 ;
        RECT 1424.350 0.690 1429.490 4.280 ;
        RECT 1430.330 0.690 1435.470 4.280 ;
        RECT 1436.310 0.690 1441.450 4.280 ;
        RECT 1442.290 0.690 1447.430 4.280 ;
        RECT 1448.270 0.690 1453.410 4.280 ;
        RECT 1454.250 0.690 1459.390 4.280 ;
        RECT 1460.230 0.690 1465.370 4.280 ;
        RECT 1466.210 0.690 1471.350 4.280 ;
        RECT 1472.190 0.690 1477.330 4.280 ;
        RECT 1478.170 0.690 1483.310 4.280 ;
        RECT 1484.150 0.690 1489.290 4.280 ;
        RECT 1490.130 0.690 1495.270 4.280 ;
        RECT 1496.110 0.690 1501.250 4.280 ;
        RECT 1502.090 0.690 1507.230 4.280 ;
        RECT 1508.070 0.690 1513.210 4.280 ;
        RECT 1514.050 0.690 1519.190 4.280 ;
        RECT 1520.030 0.690 1525.170 4.280 ;
        RECT 1526.010 0.690 1531.150 4.280 ;
        RECT 1531.990 0.690 1537.130 4.280 ;
        RECT 1537.970 0.690 1543.110 4.280 ;
        RECT 1543.950 0.690 1549.090 4.280 ;
        RECT 1549.930 0.690 1555.070 4.280 ;
        RECT 1555.910 0.690 1561.050 4.280 ;
        RECT 1561.890 0.690 1567.030 4.280 ;
        RECT 1567.870 0.690 1573.010 4.280 ;
        RECT 1573.850 0.690 1578.990 4.280 ;
        RECT 1579.830 0.690 1584.970 4.280 ;
        RECT 1585.810 0.690 1590.950 4.280 ;
        RECT 1591.790 0.690 1596.930 4.280 ;
        RECT 1597.770 0.690 1602.910 4.280 ;
        RECT 1603.750 0.690 1608.890 4.280 ;
        RECT 1609.730 0.690 1614.870 4.280 ;
        RECT 1615.710 0.690 1620.850 4.280 ;
        RECT 1621.690 0.690 1626.830 4.280 ;
        RECT 1627.670 0.690 1632.810 4.280 ;
        RECT 1633.650 0.690 1638.790 4.280 ;
        RECT 1639.630 0.690 1644.770 4.280 ;
        RECT 1645.610 0.690 1650.750 4.280 ;
        RECT 1651.590 0.690 1656.730 4.280 ;
        RECT 1657.570 0.690 1662.710 4.280 ;
        RECT 1663.550 0.690 1668.690 4.280 ;
        RECT 1669.530 0.690 1674.670 4.280 ;
        RECT 1675.510 0.690 1680.650 4.280 ;
        RECT 1681.490 0.690 1686.630 4.280 ;
        RECT 1687.470 0.690 1692.610 4.280 ;
        RECT 1693.450 0.690 1698.590 4.280 ;
        RECT 1699.430 0.690 1704.570 4.280 ;
        RECT 1705.410 0.690 1710.550 4.280 ;
        RECT 1711.390 0.690 1716.530 4.280 ;
        RECT 1717.370 0.690 1722.510 4.280 ;
        RECT 1723.350 0.690 1728.490 4.280 ;
        RECT 1729.330 0.690 1734.470 4.280 ;
        RECT 1735.310 0.690 1740.450 4.280 ;
        RECT 1741.290 0.690 1746.430 4.280 ;
        RECT 1747.270 0.690 1752.410 4.280 ;
        RECT 1753.250 0.690 1758.390 4.280 ;
        RECT 1759.230 0.690 1764.370 4.280 ;
        RECT 1765.210 0.690 1770.350 4.280 ;
        RECT 1771.190 0.690 1776.330 4.280 ;
        RECT 1777.170 0.690 1782.310 4.280 ;
        RECT 1783.150 0.690 1788.290 4.280 ;
        RECT 1789.130 0.690 1794.270 4.280 ;
        RECT 1795.110 0.690 1800.250 4.280 ;
        RECT 1801.090 0.690 1806.230 4.280 ;
        RECT 1807.070 0.690 1812.210 4.280 ;
        RECT 1813.050 0.690 1818.190 4.280 ;
        RECT 1819.030 0.690 1824.170 4.280 ;
        RECT 1825.010 0.690 1830.150 4.280 ;
        RECT 1830.990 0.690 1836.130 4.280 ;
        RECT 1836.970 0.690 1842.110 4.280 ;
        RECT 1842.950 0.690 1848.090 4.280 ;
        RECT 1848.930 0.690 1854.070 4.280 ;
        RECT 1854.910 0.690 1860.050 4.280 ;
        RECT 1860.890 0.690 1866.030 4.280 ;
        RECT 1866.870 0.690 1872.010 4.280 ;
        RECT 1872.850 0.690 1877.990 4.280 ;
        RECT 1878.830 0.690 1883.970 4.280 ;
        RECT 1884.810 0.690 1889.950 4.280 ;
        RECT 1890.790 0.690 1895.930 4.280 ;
        RECT 1896.770 0.690 1901.910 4.280 ;
        RECT 1902.750 0.690 1907.890 4.280 ;
        RECT 1908.730 0.690 1913.870 4.280 ;
        RECT 1914.710 0.690 1919.850 4.280 ;
        RECT 1920.690 0.690 1925.830 4.280 ;
        RECT 1926.670 0.690 1931.810 4.280 ;
        RECT 1932.650 0.690 1937.790 4.280 ;
        RECT 1938.630 0.690 1943.770 4.280 ;
        RECT 1944.610 0.690 1949.750 4.280 ;
        RECT 1950.590 0.690 1955.730 4.280 ;
        RECT 1956.570 0.690 1961.710 4.280 ;
        RECT 1962.550 0.690 1967.690 4.280 ;
        RECT 1968.530 0.690 1973.670 4.280 ;
        RECT 1974.510 0.690 1979.650 4.280 ;
        RECT 1980.490 0.690 1985.630 4.280 ;
        RECT 1986.470 0.690 1991.610 4.280 ;
        RECT 1992.450 0.690 1997.590 4.280 ;
        RECT 1998.430 0.690 2003.570 4.280 ;
        RECT 2004.410 0.690 2009.550 4.280 ;
        RECT 2010.390 0.690 2015.530 4.280 ;
        RECT 2016.370 0.690 2021.510 4.280 ;
        RECT 2022.350 0.690 2027.490 4.280 ;
        RECT 2028.330 0.690 2033.470 4.280 ;
        RECT 2034.310 0.690 2039.450 4.280 ;
        RECT 2040.290 0.690 2045.430 4.280 ;
        RECT 2046.270 0.690 2051.410 4.280 ;
        RECT 2052.250 0.690 2057.390 4.280 ;
        RECT 2058.230 0.690 2063.370 4.280 ;
        RECT 2064.210 0.690 2069.350 4.280 ;
        RECT 2070.190 0.690 2075.330 4.280 ;
        RECT 2076.170 0.690 2081.310 4.280 ;
        RECT 2082.150 0.690 2087.290 4.280 ;
        RECT 2088.130 0.690 2093.270 4.280 ;
        RECT 2094.110 0.690 2099.250 4.280 ;
        RECT 2100.090 0.690 2105.230 4.280 ;
        RECT 2106.070 0.690 2111.210 4.280 ;
        RECT 2112.050 0.690 2117.190 4.280 ;
        RECT 2118.030 0.690 2123.170 4.280 ;
        RECT 2124.010 0.690 2129.150 4.280 ;
        RECT 2129.990 0.690 2135.130 4.280 ;
        RECT 2135.970 0.690 2141.110 4.280 ;
        RECT 2141.950 0.690 2147.090 4.280 ;
        RECT 2147.930 0.690 2153.070 4.280 ;
        RECT 2153.910 0.690 2159.050 4.280 ;
        RECT 2159.890 0.690 2165.030 4.280 ;
        RECT 2165.870 0.690 2171.010 4.280 ;
        RECT 2171.850 0.690 2176.990 4.280 ;
        RECT 2177.830 0.690 2182.970 4.280 ;
        RECT 2183.810 0.690 2188.950 4.280 ;
        RECT 2189.790 0.690 2194.930 4.280 ;
        RECT 2195.770 0.690 2200.910 4.280 ;
        RECT 2201.750 0.690 2206.890 4.280 ;
        RECT 2207.730 0.690 2212.870 4.280 ;
        RECT 2213.710 0.690 2218.850 4.280 ;
        RECT 2219.690 0.690 2224.830 4.280 ;
        RECT 2225.670 0.690 2230.810 4.280 ;
        RECT 2231.650 0.690 2236.790 4.280 ;
        RECT 2237.630 0.690 2242.770 4.280 ;
        RECT 2243.610 0.690 2248.750 4.280 ;
        RECT 2249.590 0.690 2254.730 4.280 ;
        RECT 2255.570 0.690 2260.710 4.280 ;
        RECT 2261.550 0.690 2266.690 4.280 ;
        RECT 2267.530 0.690 2272.670 4.280 ;
        RECT 2273.510 0.690 2278.650 4.280 ;
        RECT 2279.490 0.690 2284.630 4.280 ;
        RECT 2285.470 0.690 2290.610 4.280 ;
        RECT 2291.450 0.690 2296.590 4.280 ;
        RECT 2297.430 0.690 2302.570 4.280 ;
        RECT 2303.410 0.690 2308.550 4.280 ;
        RECT 2309.390 0.690 2314.530 4.280 ;
        RECT 2315.370 0.690 2320.510 4.280 ;
        RECT 2321.350 0.690 2326.490 4.280 ;
        RECT 2327.330 0.690 2332.470 4.280 ;
        RECT 2333.310 0.690 2338.450 4.280 ;
        RECT 2339.290 0.690 2344.430 4.280 ;
        RECT 2345.270 0.690 2350.410 4.280 ;
        RECT 2351.250 0.690 2356.390 4.280 ;
        RECT 2357.230 0.690 2362.370 4.280 ;
        RECT 2363.210 0.690 2368.350 4.280 ;
        RECT 2369.190 0.690 2374.330 4.280 ;
        RECT 2375.170 0.690 2380.310 4.280 ;
        RECT 2381.150 0.690 2386.290 4.280 ;
        RECT 2387.130 0.690 2392.270 4.280 ;
        RECT 2393.110 0.690 2398.250 4.280 ;
        RECT 2399.090 0.690 2404.230 4.280 ;
        RECT 2405.070 0.690 2410.210 4.280 ;
        RECT 2411.050 0.690 2416.190 4.280 ;
        RECT 2417.030 0.690 2422.170 4.280 ;
        RECT 2423.010 0.690 2428.150 4.280 ;
        RECT 2428.990 0.690 2434.130 4.280 ;
        RECT 2434.970 0.690 2440.110 4.280 ;
        RECT 2440.950 0.690 2446.090 4.280 ;
        RECT 2446.930 0.690 2452.070 4.280 ;
        RECT 2452.910 0.690 2458.050 4.280 ;
        RECT 2458.890 0.690 2464.030 4.280 ;
        RECT 2464.870 0.690 2470.010 4.280 ;
        RECT 2470.850 0.690 2475.990 4.280 ;
        RECT 2476.830 0.690 2481.970 4.280 ;
        RECT 2482.810 0.690 2487.950 4.280 ;
        RECT 2488.790 0.690 2493.930 4.280 ;
        RECT 2494.770 0.690 2499.910 4.280 ;
        RECT 2500.750 0.690 2505.890 4.280 ;
        RECT 2506.730 0.690 2511.870 4.280 ;
        RECT 2512.710 0.690 2517.850 4.280 ;
        RECT 2518.690 0.690 2523.830 4.280 ;
        RECT 2524.670 0.690 2529.810 4.280 ;
        RECT 2530.650 0.690 2535.790 4.280 ;
        RECT 2536.630 0.690 2541.770 4.280 ;
        RECT 2542.610 0.690 2547.750 4.280 ;
        RECT 2548.590 0.690 2553.730 4.280 ;
        RECT 2554.570 0.690 2559.710 4.280 ;
        RECT 2560.550 0.690 2565.690 4.280 ;
        RECT 2566.530 0.690 2571.670 4.280 ;
        RECT 2572.510 0.690 2577.650 4.280 ;
        RECT 2578.490 0.690 2583.630 4.280 ;
        RECT 2584.470 0.690 2589.610 4.280 ;
        RECT 2590.450 0.690 2595.590 4.280 ;
        RECT 2596.430 0.690 2601.570 4.280 ;
        RECT 2602.410 0.690 2607.550 4.280 ;
        RECT 2608.390 0.690 2613.530 4.280 ;
        RECT 2614.370 0.690 2619.510 4.280 ;
        RECT 2620.350 0.690 2625.490 4.280 ;
        RECT 2626.330 0.690 2631.470 4.280 ;
        RECT 2632.310 0.690 2637.450 4.280 ;
        RECT 2638.290 0.690 2643.430 4.280 ;
        RECT 2644.270 0.690 2649.410 4.280 ;
        RECT 2650.250 0.690 2655.390 4.280 ;
        RECT 2656.230 0.690 2661.370 4.280 ;
        RECT 2662.210 0.690 2667.350 4.280 ;
        RECT 2668.190 0.690 2673.330 4.280 ;
        RECT 2674.170 0.690 2679.310 4.280 ;
        RECT 2680.150 0.690 2685.290 4.280 ;
        RECT 2686.130 0.690 2691.270 4.280 ;
        RECT 2692.110 0.690 2697.250 4.280 ;
        RECT 2698.090 0.690 2703.230 4.280 ;
        RECT 2704.070 0.690 2709.210 4.280 ;
        RECT 2710.050 0.690 2715.190 4.280 ;
        RECT 2716.030 0.690 2721.170 4.280 ;
        RECT 2722.010 0.690 2727.150 4.280 ;
        RECT 2727.990 0.690 2733.130 4.280 ;
        RECT 2733.970 0.690 2739.110 4.280 ;
        RECT 2739.950 0.690 2745.090 4.280 ;
        RECT 2745.930 0.690 2751.070 4.280 ;
        RECT 2751.910 0.690 2757.050 4.280 ;
        RECT 2757.890 0.690 2763.030 4.280 ;
        RECT 2763.870 0.690 2769.010 4.280 ;
        RECT 2769.850 0.690 2792.560 4.280 ;
      LAYER met3 ;
        RECT 4.000 2475.560 2796.000 2495.425 ;
        RECT 4.400 2474.160 2796.000 2475.560 ;
        RECT 4.000 2470.120 2796.000 2474.160 ;
        RECT 4.000 2468.720 2795.600 2470.120 ;
        RECT 4.000 2429.320 2796.000 2468.720 ;
        RECT 4.400 2427.920 2796.000 2429.320 ;
        RECT 4.000 2423.200 2796.000 2427.920 ;
        RECT 4.000 2421.800 2795.600 2423.200 ;
        RECT 4.000 2383.080 2796.000 2421.800 ;
        RECT 4.400 2381.680 2796.000 2383.080 ;
        RECT 4.000 2376.280 2796.000 2381.680 ;
        RECT 4.000 2374.880 2795.600 2376.280 ;
        RECT 4.000 2336.840 2796.000 2374.880 ;
        RECT 4.400 2335.440 2796.000 2336.840 ;
        RECT 4.000 2329.360 2796.000 2335.440 ;
        RECT 4.000 2327.960 2795.600 2329.360 ;
        RECT 4.000 2290.600 2796.000 2327.960 ;
        RECT 4.400 2289.200 2796.000 2290.600 ;
        RECT 4.000 2282.440 2796.000 2289.200 ;
        RECT 4.000 2281.040 2795.600 2282.440 ;
        RECT 4.000 2244.360 2796.000 2281.040 ;
        RECT 4.400 2242.960 2796.000 2244.360 ;
        RECT 4.000 2235.520 2796.000 2242.960 ;
        RECT 4.000 2234.120 2795.600 2235.520 ;
        RECT 4.000 2198.120 2796.000 2234.120 ;
        RECT 4.400 2196.720 2796.000 2198.120 ;
        RECT 4.000 2188.600 2796.000 2196.720 ;
        RECT 4.000 2187.200 2795.600 2188.600 ;
        RECT 4.000 2151.880 2796.000 2187.200 ;
        RECT 4.400 2150.480 2796.000 2151.880 ;
        RECT 4.000 2141.680 2796.000 2150.480 ;
        RECT 4.000 2140.280 2795.600 2141.680 ;
        RECT 4.000 2105.640 2796.000 2140.280 ;
        RECT 4.400 2104.240 2796.000 2105.640 ;
        RECT 4.000 2094.760 2796.000 2104.240 ;
        RECT 4.000 2093.360 2795.600 2094.760 ;
        RECT 4.000 2059.400 2796.000 2093.360 ;
        RECT 4.400 2058.000 2796.000 2059.400 ;
        RECT 4.000 2047.840 2796.000 2058.000 ;
        RECT 4.000 2046.440 2795.600 2047.840 ;
        RECT 4.000 2013.160 2796.000 2046.440 ;
        RECT 4.400 2011.760 2796.000 2013.160 ;
        RECT 4.000 2000.920 2796.000 2011.760 ;
        RECT 4.000 1999.520 2795.600 2000.920 ;
        RECT 4.000 1966.920 2796.000 1999.520 ;
        RECT 4.400 1965.520 2796.000 1966.920 ;
        RECT 4.000 1954.000 2796.000 1965.520 ;
        RECT 4.000 1952.600 2795.600 1954.000 ;
        RECT 4.000 1920.680 2796.000 1952.600 ;
        RECT 4.400 1919.280 2796.000 1920.680 ;
        RECT 4.000 1907.080 2796.000 1919.280 ;
        RECT 4.000 1905.680 2795.600 1907.080 ;
        RECT 4.000 1874.440 2796.000 1905.680 ;
        RECT 4.400 1873.040 2796.000 1874.440 ;
        RECT 4.000 1860.160 2796.000 1873.040 ;
        RECT 4.000 1858.760 2795.600 1860.160 ;
        RECT 4.000 1828.200 2796.000 1858.760 ;
        RECT 4.400 1826.800 2796.000 1828.200 ;
        RECT 4.000 1813.240 2796.000 1826.800 ;
        RECT 4.000 1811.840 2795.600 1813.240 ;
        RECT 4.000 1781.960 2796.000 1811.840 ;
        RECT 4.400 1780.560 2796.000 1781.960 ;
        RECT 4.000 1766.320 2796.000 1780.560 ;
        RECT 4.000 1764.920 2795.600 1766.320 ;
        RECT 4.000 1735.720 2796.000 1764.920 ;
        RECT 4.400 1734.320 2796.000 1735.720 ;
        RECT 4.000 1719.400 2796.000 1734.320 ;
        RECT 4.000 1718.000 2795.600 1719.400 ;
        RECT 4.000 1689.480 2796.000 1718.000 ;
        RECT 4.400 1688.080 2796.000 1689.480 ;
        RECT 4.000 1672.480 2796.000 1688.080 ;
        RECT 4.000 1671.080 2795.600 1672.480 ;
        RECT 4.000 1643.240 2796.000 1671.080 ;
        RECT 4.400 1641.840 2796.000 1643.240 ;
        RECT 4.000 1625.560 2796.000 1641.840 ;
        RECT 4.000 1624.160 2795.600 1625.560 ;
        RECT 4.000 1597.000 2796.000 1624.160 ;
        RECT 4.400 1595.600 2796.000 1597.000 ;
        RECT 4.000 1578.640 2796.000 1595.600 ;
        RECT 4.000 1577.240 2795.600 1578.640 ;
        RECT 4.000 1550.760 2796.000 1577.240 ;
        RECT 4.400 1549.360 2796.000 1550.760 ;
        RECT 4.000 1531.720 2796.000 1549.360 ;
        RECT 4.000 1530.320 2795.600 1531.720 ;
        RECT 4.000 1504.520 2796.000 1530.320 ;
        RECT 4.400 1503.120 2796.000 1504.520 ;
        RECT 4.000 1484.800 2796.000 1503.120 ;
        RECT 4.000 1483.400 2795.600 1484.800 ;
        RECT 4.000 1458.280 2796.000 1483.400 ;
        RECT 4.400 1456.880 2796.000 1458.280 ;
        RECT 4.000 1437.880 2796.000 1456.880 ;
        RECT 4.000 1436.480 2795.600 1437.880 ;
        RECT 4.000 1412.040 2796.000 1436.480 ;
        RECT 4.400 1410.640 2796.000 1412.040 ;
        RECT 4.000 1390.960 2796.000 1410.640 ;
        RECT 4.000 1389.560 2795.600 1390.960 ;
        RECT 4.000 1365.800 2796.000 1389.560 ;
        RECT 4.400 1364.400 2796.000 1365.800 ;
        RECT 4.000 1344.040 2796.000 1364.400 ;
        RECT 4.000 1342.640 2795.600 1344.040 ;
        RECT 4.000 1319.560 2796.000 1342.640 ;
        RECT 4.400 1318.160 2796.000 1319.560 ;
        RECT 4.000 1297.120 2796.000 1318.160 ;
        RECT 4.000 1295.720 2795.600 1297.120 ;
        RECT 4.000 1273.320 2796.000 1295.720 ;
        RECT 4.400 1271.920 2796.000 1273.320 ;
        RECT 4.000 1250.200 2796.000 1271.920 ;
        RECT 4.000 1248.800 2795.600 1250.200 ;
        RECT 4.000 1227.080 2796.000 1248.800 ;
        RECT 4.400 1225.680 2796.000 1227.080 ;
        RECT 4.000 1203.280 2796.000 1225.680 ;
        RECT 4.000 1201.880 2795.600 1203.280 ;
        RECT 4.000 1180.840 2796.000 1201.880 ;
        RECT 4.400 1179.440 2796.000 1180.840 ;
        RECT 4.000 1156.360 2796.000 1179.440 ;
        RECT 4.000 1154.960 2795.600 1156.360 ;
        RECT 4.000 1134.600 2796.000 1154.960 ;
        RECT 4.400 1133.200 2796.000 1134.600 ;
        RECT 4.000 1109.440 2796.000 1133.200 ;
        RECT 4.000 1108.040 2795.600 1109.440 ;
        RECT 4.000 1088.360 2796.000 1108.040 ;
        RECT 4.400 1086.960 2796.000 1088.360 ;
        RECT 4.000 1062.520 2796.000 1086.960 ;
        RECT 4.000 1061.120 2795.600 1062.520 ;
        RECT 4.000 1042.120 2796.000 1061.120 ;
        RECT 4.400 1040.720 2796.000 1042.120 ;
        RECT 4.000 1015.600 2796.000 1040.720 ;
        RECT 4.000 1014.200 2795.600 1015.600 ;
        RECT 4.000 995.880 2796.000 1014.200 ;
        RECT 4.400 994.480 2796.000 995.880 ;
        RECT 4.000 968.680 2796.000 994.480 ;
        RECT 4.000 967.280 2795.600 968.680 ;
        RECT 4.000 949.640 2796.000 967.280 ;
        RECT 4.400 948.240 2796.000 949.640 ;
        RECT 4.000 921.760 2796.000 948.240 ;
        RECT 4.000 920.360 2795.600 921.760 ;
        RECT 4.000 903.400 2796.000 920.360 ;
        RECT 4.400 902.000 2796.000 903.400 ;
        RECT 4.000 874.840 2796.000 902.000 ;
        RECT 4.000 873.440 2795.600 874.840 ;
        RECT 4.000 857.160 2796.000 873.440 ;
        RECT 4.400 855.760 2796.000 857.160 ;
        RECT 4.000 827.920 2796.000 855.760 ;
        RECT 4.000 826.520 2795.600 827.920 ;
        RECT 4.000 810.920 2796.000 826.520 ;
        RECT 4.400 809.520 2796.000 810.920 ;
        RECT 4.000 781.000 2796.000 809.520 ;
        RECT 4.000 779.600 2795.600 781.000 ;
        RECT 4.000 764.680 2796.000 779.600 ;
        RECT 4.400 763.280 2796.000 764.680 ;
        RECT 4.000 734.080 2796.000 763.280 ;
        RECT 4.000 732.680 2795.600 734.080 ;
        RECT 4.000 718.440 2796.000 732.680 ;
        RECT 4.400 717.040 2796.000 718.440 ;
        RECT 4.000 687.160 2796.000 717.040 ;
        RECT 4.000 685.760 2795.600 687.160 ;
        RECT 4.000 672.200 2796.000 685.760 ;
        RECT 4.400 670.800 2796.000 672.200 ;
        RECT 4.000 640.240 2796.000 670.800 ;
        RECT 4.000 638.840 2795.600 640.240 ;
        RECT 4.000 625.960 2796.000 638.840 ;
        RECT 4.400 624.560 2796.000 625.960 ;
        RECT 4.000 593.320 2796.000 624.560 ;
        RECT 4.000 591.920 2795.600 593.320 ;
        RECT 4.000 579.720 2796.000 591.920 ;
        RECT 4.400 578.320 2796.000 579.720 ;
        RECT 4.000 546.400 2796.000 578.320 ;
        RECT 4.000 545.000 2795.600 546.400 ;
        RECT 4.000 533.480 2796.000 545.000 ;
        RECT 4.400 532.080 2796.000 533.480 ;
        RECT 4.000 499.480 2796.000 532.080 ;
        RECT 4.000 498.080 2795.600 499.480 ;
        RECT 4.000 487.240 2796.000 498.080 ;
        RECT 4.400 485.840 2796.000 487.240 ;
        RECT 4.000 452.560 2796.000 485.840 ;
        RECT 4.000 451.160 2795.600 452.560 ;
        RECT 4.000 441.000 2796.000 451.160 ;
        RECT 4.400 439.600 2796.000 441.000 ;
        RECT 4.000 405.640 2796.000 439.600 ;
        RECT 4.000 404.240 2795.600 405.640 ;
        RECT 4.000 394.760 2796.000 404.240 ;
        RECT 4.400 393.360 2796.000 394.760 ;
        RECT 4.000 358.720 2796.000 393.360 ;
        RECT 4.000 357.320 2795.600 358.720 ;
        RECT 4.000 348.520 2796.000 357.320 ;
        RECT 4.400 347.120 2796.000 348.520 ;
        RECT 4.000 311.800 2796.000 347.120 ;
        RECT 4.000 310.400 2795.600 311.800 ;
        RECT 4.000 302.280 2796.000 310.400 ;
        RECT 4.400 300.880 2796.000 302.280 ;
        RECT 4.000 264.880 2796.000 300.880 ;
        RECT 4.000 263.480 2795.600 264.880 ;
        RECT 4.000 256.040 2796.000 263.480 ;
        RECT 4.400 254.640 2796.000 256.040 ;
        RECT 4.000 217.960 2796.000 254.640 ;
        RECT 4.000 216.560 2795.600 217.960 ;
        RECT 4.000 209.800 2796.000 216.560 ;
        RECT 4.400 208.400 2796.000 209.800 ;
        RECT 4.000 171.040 2796.000 208.400 ;
        RECT 4.000 169.640 2795.600 171.040 ;
        RECT 4.000 163.560 2796.000 169.640 ;
        RECT 4.400 162.160 2796.000 163.560 ;
        RECT 4.000 124.120 2796.000 162.160 ;
        RECT 4.000 122.720 2795.600 124.120 ;
        RECT 4.000 117.320 2796.000 122.720 ;
        RECT 4.400 115.920 2796.000 117.320 ;
        RECT 4.000 77.200 2796.000 115.920 ;
        RECT 4.000 75.800 2795.600 77.200 ;
        RECT 4.000 71.080 2796.000 75.800 ;
        RECT 4.400 69.680 2796.000 71.080 ;
        RECT 4.000 30.280 2796.000 69.680 ;
        RECT 4.000 28.880 2795.600 30.280 ;
        RECT 4.000 24.840 2796.000 28.880 ;
        RECT 4.400 23.440 2796.000 24.840 ;
        RECT 4.000 2.215 2796.000 23.440 ;
      LAYER met4 ;
        RECT 87.695 2489.440 2731.185 2495.425 ;
        RECT 87.695 10.240 97.440 2489.440 ;
        RECT 99.840 10.240 174.240 2489.440 ;
        RECT 176.640 10.240 251.040 2489.440 ;
        RECT 253.440 10.240 327.840 2489.440 ;
        RECT 330.240 10.240 404.640 2489.440 ;
        RECT 407.040 10.240 481.440 2489.440 ;
        RECT 483.840 10.240 558.240 2489.440 ;
        RECT 560.640 10.240 635.040 2489.440 ;
        RECT 637.440 10.240 711.840 2489.440 ;
        RECT 714.240 10.240 788.640 2489.440 ;
        RECT 791.040 10.240 865.440 2489.440 ;
        RECT 867.840 10.240 942.240 2489.440 ;
        RECT 944.640 10.240 1019.040 2489.440 ;
        RECT 1021.440 10.240 1095.840 2489.440 ;
        RECT 1098.240 10.240 1172.640 2489.440 ;
        RECT 1175.040 10.240 1249.440 2489.440 ;
        RECT 1251.840 10.240 1326.240 2489.440 ;
        RECT 1328.640 10.240 1403.040 2489.440 ;
        RECT 1405.440 10.240 1479.840 2489.440 ;
        RECT 1482.240 10.240 1556.640 2489.440 ;
        RECT 1559.040 10.240 1633.440 2489.440 ;
        RECT 1635.840 10.240 1710.240 2489.440 ;
        RECT 1712.640 10.240 1787.040 2489.440 ;
        RECT 1789.440 10.240 1863.840 2489.440 ;
        RECT 1866.240 10.240 1940.640 2489.440 ;
        RECT 1943.040 10.240 2017.440 2489.440 ;
        RECT 2019.840 10.240 2094.240 2489.440 ;
        RECT 2096.640 10.240 2171.040 2489.440 ;
        RECT 2173.440 10.240 2247.840 2489.440 ;
        RECT 2250.240 10.240 2324.640 2489.440 ;
        RECT 2327.040 10.240 2401.440 2489.440 ;
        RECT 2403.840 10.240 2478.240 2489.440 ;
        RECT 2480.640 10.240 2555.040 2489.440 ;
        RECT 2557.440 10.240 2631.840 2489.440 ;
        RECT 2634.240 10.240 2708.640 2489.440 ;
        RECT 2711.040 10.240 2731.185 2489.440 ;
        RECT 87.695 2.895 2731.185 10.240 ;
  END
END soomrv
END LIBRARY

